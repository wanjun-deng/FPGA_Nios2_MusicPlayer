// mysystem.v

// Generated using ACDS version 13.0 156 at 2025.12.27.21:41:46

`timescale 1 ps / 1 ps
module mysystem (
		input  wire       clk_clk,                     //               clk.clk
		input  wire       reset_reset_n,               //             reset.reset_n
		output wire [7:0] led_export,                  //               led.export
		output wire       vib_export_export,           //        vib_export.export
		input  wire [3:0] keyboard_export_Row_i,       //   keyboard_export.Row_i
		output wire [3:0] keyboard_export_Col_o,       //                  .Col_o
		input  wire       ir_decode_export_iIR,        //  ir_decode_export.iIR
		output wire       ir_decode_export_Get_Flag_o, //                  .Get_Flag_o
		output wire       hex_driver_export_SH_CP,     // hex_driver_export.SH_CP
		output wire       hex_driver_export_ST_CP,     //                  .ST_CP
		output wire       hex_driver_export_DS         //                  .DS
	);

	wire         nios2_instruction_master_waitrequest;                                                                // nios2_instruction_master_translator:av_waitrequest -> nios2:i_waitrequest
	wire  [15:0] nios2_instruction_master_address;                                                                    // nios2:i_address -> nios2_instruction_master_translator:av_address
	wire         nios2_instruction_master_read;                                                                       // nios2:i_read -> nios2_instruction_master_translator:av_read
	wire  [31:0] nios2_instruction_master_readdata;                                                                   // nios2_instruction_master_translator:av_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_readdatavalid;                                                              // nios2_instruction_master_translator:av_readdatavalid -> nios2:i_readdatavalid
	wire         nios2_data_master_waitrequest;                                                                       // nios2_data_master_translator:av_waitrequest -> nios2:d_waitrequest
	wire  [31:0] nios2_data_master_writedata;                                                                         // nios2:d_writedata -> nios2_data_master_translator:av_writedata
	wire  [15:0] nios2_data_master_address;                                                                           // nios2:d_address -> nios2_data_master_translator:av_address
	wire         nios2_data_master_write;                                                                             // nios2:d_write -> nios2_data_master_translator:av_write
	wire         nios2_data_master_read;                                                                              // nios2:d_read -> nios2_data_master_translator:av_read
	wire  [31:0] nios2_data_master_readdata;                                                                          // nios2_data_master_translator:av_readdata -> nios2:d_readdata
	wire         nios2_data_master_debugaccess;                                                                       // nios2:jtag_debug_module_debugaccess_to_roms -> nios2_data_master_translator:av_debugaccess
	wire         nios2_data_master_readdatavalid;                                                                     // nios2_data_master_translator:av_readdatavalid -> nios2:d_readdatavalid
	wire   [3:0] nios2_data_master_byteenable;                                                                        // nios2:d_byteenable -> nios2_data_master_translator:av_byteenable
	wire         nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                  // nios2:jtag_debug_module_waitrequest -> nios2_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                    // nios2_jtag_debug_module_translator:av_writedata -> nios2:jtag_debug_module_writedata
	wire   [8:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_address;                                      // nios2_jtag_debug_module_translator:av_address -> nios2:jtag_debug_module_address
	wire         nios2_jtag_debug_module_translator_avalon_anti_slave_0_write;                                        // nios2_jtag_debug_module_translator:av_write -> nios2:jtag_debug_module_write
	wire         nios2_jtag_debug_module_translator_avalon_anti_slave_0_read;                                         // nios2_jtag_debug_module_translator:av_read -> nios2:jtag_debug_module_read
	wire  [31:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                     // nios2:jtag_debug_module_readdata -> nios2_jtag_debug_module_translator:av_readdata
	wire         nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                  // nios2_jtag_debug_module_translator:av_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [3:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                   // nios2_jtag_debug_module_translator:av_byteenable -> nios2:jtag_debug_module_byteenable
	wire  [31:0] rom_s1_translator_avalon_anti_slave_0_writedata;                                                     // rom_s1_translator:av_writedata -> rom:writedata
	wire   [8:0] rom_s1_translator_avalon_anti_slave_0_address;                                                       // rom_s1_translator:av_address -> rom:address
	wire         rom_s1_translator_avalon_anti_slave_0_chipselect;                                                    // rom_s1_translator:av_chipselect -> rom:chipselect
	wire         rom_s1_translator_avalon_anti_slave_0_clken;                                                         // rom_s1_translator:av_clken -> rom:clken
	wire         rom_s1_translator_avalon_anti_slave_0_write;                                                         // rom_s1_translator:av_write -> rom:write
	wire  [31:0] rom_s1_translator_avalon_anti_slave_0_readdata;                                                      // rom:readdata -> rom_s1_translator:av_readdata
	wire         rom_s1_translator_avalon_anti_slave_0_debugaccess;                                                   // rom_s1_translator:av_debugaccess -> rom:debugaccess
	wire   [3:0] rom_s1_translator_avalon_anti_slave_0_byteenable;                                                    // rom_s1_translator:av_byteenable -> rom:byteenable
	wire  [31:0] ram_s1_translator_avalon_anti_slave_0_writedata;                                                     // ram_s1_translator:av_writedata -> ram:writedata
	wire  [11:0] ram_s1_translator_avalon_anti_slave_0_address;                                                       // ram_s1_translator:av_address -> ram:address
	wire         ram_s1_translator_avalon_anti_slave_0_chipselect;                                                    // ram_s1_translator:av_chipselect -> ram:chipselect
	wire         ram_s1_translator_avalon_anti_slave_0_clken;                                                         // ram_s1_translator:av_clken -> ram:clken
	wire         ram_s1_translator_avalon_anti_slave_0_write;                                                         // ram_s1_translator:av_write -> ram:write
	wire  [31:0] ram_s1_translator_avalon_anti_slave_0_readdata;                                                      // ram:readdata -> ram_s1_translator:av_readdata
	wire   [3:0] ram_s1_translator_avalon_anti_slave_0_byteenable;                                                    // ram_s1_translator:av_byteenable -> ram:byteenable
	wire   [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                          // sysid_control_slave_translator:av_address -> sysid:address
	wire  [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                         // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire  [31:0] pio_led_s1_translator_avalon_anti_slave_0_writedata;                                                 // pio_led_s1_translator:av_writedata -> pio_led:writedata
	wire   [2:0] pio_led_s1_translator_avalon_anti_slave_0_address;                                                   // pio_led_s1_translator:av_address -> pio_led:address
	wire         pio_led_s1_translator_avalon_anti_slave_0_chipselect;                                                // pio_led_s1_translator:av_chipselect -> pio_led:chipselect
	wire         pio_led_s1_translator_avalon_anti_slave_0_write;                                                     // pio_led_s1_translator:av_write -> pio_led:write_n
	wire  [31:0] pio_led_s1_translator_avalon_anti_slave_0_readdata;                                                  // pio_led:readdata -> pio_led_s1_translator:av_readdata
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                 // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire   [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                   // timer_0_s1_translator:av_address -> timer_0:address
	wire         timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                                // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire         timer_0_s1_translator_avalon_anti_slave_0_write;                                                     // timer_0_s1_translator:av_write -> timer_0:write_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                  // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                            // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                              // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                             // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                   // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                               // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire   [7:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                              // FreqSynth_IP_0_avalon_slave_0_translator:av_writedata -> FreqSynth_IP_0:writedata
	wire   [1:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                // FreqSynth_IP_0_avalon_slave_0_translator:av_address -> FreqSynth_IP_0:address
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                             // FreqSynth_IP_0_avalon_slave_0_translator:av_chipselect -> FreqSynth_IP_0:chipselect
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                  // FreqSynth_IP_0_avalon_slave_0_translator:av_write -> FreqSynth_IP_0:write
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                   // FreqSynth_IP_0_avalon_slave_0_translator:av_read -> FreqSynth_IP_0:read
	wire   [7:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                               // FreqSynth_IP_0:readdata -> FreqSynth_IP_0_avalon_slave_0_translator:av_readdata
	wire   [7:0] keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                               // KeyBoard_IP_0_avalon_slave_0_translator:av_writedata -> KeyBoard_IP_0:writedata
	wire   [0:0] keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                 // KeyBoard_IP_0_avalon_slave_0_translator:av_address -> KeyBoard_IP_0:address
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                              // KeyBoard_IP_0_avalon_slave_0_translator:av_chipselect -> KeyBoard_IP_0:chipselect
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                   // KeyBoard_IP_0_avalon_slave_0_translator:av_write -> KeyBoard_IP_0:write
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                    // KeyBoard_IP_0_avalon_slave_0_translator:av_read -> KeyBoard_IP_0:read
	wire   [7:0] keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                // KeyBoard_IP_0:readdata -> KeyBoard_IP_0_avalon_slave_0_translator:av_readdata
	wire   [7:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                              // Ir_Decode_IP_0_avalon_slave_0_translator:av_writedata -> Ir_Decode_IP_0:writedata
	wire   [2:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                // Ir_Decode_IP_0_avalon_slave_0_translator:av_address -> Ir_Decode_IP_0:address
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                             // Ir_Decode_IP_0_avalon_slave_0_translator:av_chipselect -> Ir_Decode_IP_0:chipselect
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                  // Ir_Decode_IP_0_avalon_slave_0_translator:av_write -> Ir_Decode_IP_0:write
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                   // Ir_Decode_IP_0_avalon_slave_0_translator:av_read -> Ir_Decode_IP_0:read
	wire   [7:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                               // Ir_Decode_IP_0:readdata -> Ir_Decode_IP_0_avalon_slave_0_translator:av_readdata
	wire   [7:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                             // Hex_Driver_IP_0_avalon_slave_0_translator:av_writedata -> Hex_Driver_IP_0:writedata
	wire   [2:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                               // Hex_Driver_IP_0_avalon_slave_0_translator:av_address -> Hex_Driver_IP_0:address
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                            // Hex_Driver_IP_0_avalon_slave_0_translator:av_chipselect -> Hex_Driver_IP_0:chipselect
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                 // Hex_Driver_IP_0_avalon_slave_0_translator:av_write -> Hex_Driver_IP_0:write
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                  // Hex_Driver_IP_0_avalon_slave_0_translator:av_read -> Hex_Driver_IP_0:read
	wire   [7:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                              // Hex_Driver_IP_0:readdata -> Hex_Driver_IP_0_avalon_slave_0_translator:av_readdata
	wire         nios2_instruction_master_translator_avalon_universal_master_0_waitrequest;                           // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_instruction_master_translator_avalon_universal_master_0_burstcount;                            // nios2_instruction_master_translator:uav_burstcount -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_instruction_master_translator_avalon_universal_master_0_writedata;                             // nios2_instruction_master_translator:uav_writedata -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [15:0] nios2_instruction_master_translator_avalon_universal_master_0_address;                               // nios2_instruction_master_translator:uav_address -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_instruction_master_translator_avalon_universal_master_0_lock;                                  // nios2_instruction_master_translator:uav_lock -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_instruction_master_translator_avalon_universal_master_0_write;                                 // nios2_instruction_master_translator:uav_write -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_instruction_master_translator_avalon_universal_master_0_read;                                  // nios2_instruction_master_translator:uav_read -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_instruction_master_translator_avalon_universal_master_0_readdata;                              // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_instruction_master_translator:uav_readdata
	wire         nios2_instruction_master_translator_avalon_universal_master_0_debugaccess;                           // nios2_instruction_master_translator:uav_debugaccess -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_instruction_master_translator_avalon_universal_master_0_byteenable;                            // nios2_instruction_master_translator:uav_byteenable -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid;                         // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_instruction_master_translator:uav_readdatavalid
	wire         nios2_data_master_translator_avalon_universal_master_0_waitrequest;                                  // nios2_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_data_master_translator_avalon_universal_master_0_burstcount;                                   // nios2_data_master_translator:uav_burstcount -> nios2_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_data_master_translator_avalon_universal_master_0_writedata;                                    // nios2_data_master_translator:uav_writedata -> nios2_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [15:0] nios2_data_master_translator_avalon_universal_master_0_address;                                      // nios2_data_master_translator:uav_address -> nios2_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_data_master_translator_avalon_universal_master_0_lock;                                         // nios2_data_master_translator:uav_lock -> nios2_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_data_master_translator_avalon_universal_master_0_write;                                        // nios2_data_master_translator:uav_write -> nios2_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_data_master_translator_avalon_universal_master_0_read;                                         // nios2_data_master_translator:uav_read -> nios2_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_data_master_translator_avalon_universal_master_0_readdata;                                     // nios2_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_data_master_translator:uav_readdata
	wire         nios2_data_master_translator_avalon_universal_master_0_debugaccess;                                  // nios2_data_master_translator:uav_debugaccess -> nios2_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_data_master_translator_avalon_universal_master_0_byteenable;                                   // nios2_data_master_translator:uav_byteenable -> nios2_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_data_master_translator_avalon_universal_master_0_readdatavalid;                                // nios2_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_data_master_translator:uav_readdatavalid
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // nios2_jtag_debug_module_translator:uav_waitrequest -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                      // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_jtag_debug_module_translator:uav_writedata
	wire  [15:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                        // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_jtag_debug_module_translator:uav_address
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                          // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_jtag_debug_module_translator:uav_write
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                           // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_jtag_debug_module_translator:uav_lock
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                           // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                       // nios2_jtag_debug_module_translator:uav_readdata -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // nios2_jtag_debug_module_translator:uav_readdatavalid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_jtag_debug_module_translator:uav_byteenable
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [91:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                    // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [91:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         rom_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // rom_s1_translator:uav_waitrequest -> rom_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] rom_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // rom_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> rom_s1_translator:uav_burstcount
	wire  [31:0] rom_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // rom_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> rom_s1_translator:uav_writedata
	wire  [15:0] rom_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // rom_s1_translator_avalon_universal_slave_0_agent:m0_address -> rom_s1_translator:uav_address
	wire         rom_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // rom_s1_translator_avalon_universal_slave_0_agent:m0_write -> rom_s1_translator:uav_write
	wire         rom_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // rom_s1_translator_avalon_universal_slave_0_agent:m0_lock -> rom_s1_translator:uav_lock
	wire         rom_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // rom_s1_translator_avalon_universal_slave_0_agent:m0_read -> rom_s1_translator:uav_read
	wire  [31:0] rom_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // rom_s1_translator:uav_readdata -> rom_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         rom_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // rom_s1_translator:uav_readdatavalid -> rom_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         rom_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // rom_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> rom_s1_translator:uav_debugaccess
	wire   [3:0] rom_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // rom_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> rom_s1_translator:uav_byteenable
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // rom_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // rom_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // rom_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [91:0] rom_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // rom_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> rom_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> rom_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> rom_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> rom_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [91:0] rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> rom_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // rom_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // rom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> rom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // rom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> rom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // rom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> rom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // ram_s1_translator:uav_waitrequest -> ram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // ram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ram_s1_translator:uav_burstcount
	wire  [31:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // ram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ram_s1_translator:uav_writedata
	wire  [15:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // ram_s1_translator_avalon_universal_slave_0_agent:m0_address -> ram_s1_translator:uav_address
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // ram_s1_translator_avalon_universal_slave_0_agent:m0_write -> ram_s1_translator:uav_write
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // ram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ram_s1_translator:uav_lock
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // ram_s1_translator_avalon_universal_slave_0_agent:m0_read -> ram_s1_translator:uav_read
	wire  [31:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // ram_s1_translator:uav_readdata -> ram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // ram_s1_translator:uav_readdatavalid -> ram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // ram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ram_s1_translator:uav_debugaccess
	wire   [3:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // ram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ram_s1_translator:uav_byteenable
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // ram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // ram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // ram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [91:0] ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // ram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [91:0] ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire  [15:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [91:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [91:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // pio_led_s1_translator:uav_waitrequest -> pio_led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_led_s1_translator:uav_burstcount
	wire  [31:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_led_s1_translator:uav_writedata
	wire  [15:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_led_s1_translator:uav_address
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_led_s1_translator:uav_write
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_led_s1_translator:uav_lock
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_led_s1_translator:uav_read
	wire  [31:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // pio_led_s1_translator:uav_readdata -> pio_led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // pio_led_s1_translator:uav_readdatavalid -> pio_led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_led_s1_translator:uav_debugaccess
	wire   [3:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_led_s1_translator:uav_byteenable
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [91:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [91:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire  [15:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [91:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [91:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [15:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [91:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [91:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // FreqSynth_IP_0_avalon_slave_0_translator:uav_waitrequest -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [0:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;               // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> FreqSynth_IP_0_avalon_slave_0_translator:uav_burstcount
	wire   [7:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> FreqSynth_IP_0_avalon_slave_0_translator:uav_writedata
	wire  [15:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                  // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> FreqSynth_IP_0_avalon_slave_0_translator:uav_address
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                    // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> FreqSynth_IP_0_avalon_slave_0_translator:uav_write
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                     // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> FreqSynth_IP_0_avalon_slave_0_translator:uav_lock
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                     // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> FreqSynth_IP_0_avalon_slave_0_translator:uav_read
	wire   [7:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                 // FreqSynth_IP_0_avalon_slave_0_translator:uav_readdata -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // FreqSynth_IP_0_avalon_slave_0_translator:uav_readdatavalid -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FreqSynth_IP_0_avalon_slave_0_translator:uav_debugaccess
	wire   [0:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;               // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> FreqSynth_IP_0_avalon_slave_0_translator:uav_byteenable
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;             // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [64:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;              // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;             // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [64:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [9:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // KeyBoard_IP_0_avalon_slave_0_translator:uav_waitrequest -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [0:0] keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> KeyBoard_IP_0_avalon_slave_0_translator:uav_burstcount
	wire   [7:0] keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                 // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> KeyBoard_IP_0_avalon_slave_0_translator:uav_writedata
	wire  [15:0] keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                   // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> KeyBoard_IP_0_avalon_slave_0_translator:uav_address
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                     // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> KeyBoard_IP_0_avalon_slave_0_translator:uav_write
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                      // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> KeyBoard_IP_0_avalon_slave_0_translator:uav_lock
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                      // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> KeyBoard_IP_0_avalon_slave_0_translator:uav_read
	wire   [7:0] keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                  // KeyBoard_IP_0_avalon_slave_0_translator:uav_readdata -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // KeyBoard_IP_0_avalon_slave_0_translator:uav_readdatavalid -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> KeyBoard_IP_0_avalon_slave_0_translator:uav_debugaccess
	wire   [0:0] keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> KeyBoard_IP_0_avalon_slave_0_translator:uav_byteenable
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;              // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [64:0] keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;               // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;              // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [64:0] keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [9:0] keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Ir_Decode_IP_0_avalon_slave_0_translator:uav_waitrequest -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [0:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Ir_Decode_IP_0_avalon_slave_0_translator:uav_burstcount
	wire   [7:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Ir_Decode_IP_0_avalon_slave_0_translator:uav_writedata
	wire  [15:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                  // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Ir_Decode_IP_0_avalon_slave_0_translator:uav_address
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                    // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Ir_Decode_IP_0_avalon_slave_0_translator:uav_write
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                     // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Ir_Decode_IP_0_avalon_slave_0_translator:uav_lock
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                     // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Ir_Decode_IP_0_avalon_slave_0_translator:uav_read
	wire   [7:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Ir_Decode_IP_0_avalon_slave_0_translator:uav_readdata -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Ir_Decode_IP_0_avalon_slave_0_translator:uav_readdatavalid -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Ir_Decode_IP_0_avalon_slave_0_translator:uav_debugaccess
	wire   [0:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Ir_Decode_IP_0_avalon_slave_0_translator:uav_byteenable
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [64:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;              // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [64:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [9:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Hex_Driver_IP_0_avalon_slave_0_translator:uav_waitrequest -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [0:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Hex_Driver_IP_0_avalon_slave_0_translator:uav_burstcount
	wire   [7:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;               // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Hex_Driver_IP_0_avalon_slave_0_translator:uav_writedata
	wire  [15:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                 // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Hex_Driver_IP_0_avalon_slave_0_translator:uav_address
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                   // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Hex_Driver_IP_0_avalon_slave_0_translator:uav_write
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                    // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Hex_Driver_IP_0_avalon_slave_0_translator:uav_lock
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                    // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Hex_Driver_IP_0_avalon_slave_0_translator:uav_read
	wire   [7:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                // Hex_Driver_IP_0_avalon_slave_0_translator:uav_readdata -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Hex_Driver_IP_0_avalon_slave_0_translator:uav_readdatavalid -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Hex_Driver_IP_0_avalon_slave_0_translator:uav_debugaccess
	wire   [0:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Hex_Driver_IP_0_avalon_slave_0_translator:uav_byteenable
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [64:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;             // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [64:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [9:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                        // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [90:0] nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                         // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router:sink_ready -> nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // nios2_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid;                               // nios2_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // nios2_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [90:0] nios2_data_master_translator_avalon_universal_master_0_agent_cp_data;                                // nios2_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router_001:sink_ready -> nios2_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                          // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [90:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                           // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router:sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // rom_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // rom_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // rom_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [90:0] rom_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // rom_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         rom_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_001:sink_ready -> rom_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // ram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // ram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // ram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [90:0] ram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // ram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_002:sink_ready -> ram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [90:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_003:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [90:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         pio_led_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_004:sink_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [90:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_005:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [90:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_006:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                    // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [63:0] freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                     // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_007:sink_ready -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                     // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [63:0] keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                      // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_008:sink_ready -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                    // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [63:0] ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                     // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_009:sink_ready -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                   // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [63:0] hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                    // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_010:sink_ready -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                         // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                               // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                       // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [90:0] addr_router_src_data;                                                                                // addr_router:src_data -> limiter:cmd_sink_data
	wire  [10:0] addr_router_src_channel;                                                                             // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                               // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                         // limiter:rsp_src_endofpacket -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                               // limiter:rsp_src_valid -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                       // limiter:rsp_src_startofpacket -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [90:0] limiter_rsp_src_data;                                                                                // limiter:rsp_src_data -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [10:0] limiter_rsp_src_channel;                                                                             // limiter:rsp_src_channel -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                               // nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                     // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                           // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                   // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [90:0] addr_router_001_src_data;                                                                            // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire  [10:0] addr_router_001_src_channel;                                                                         // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                           // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                     // limiter_001:rsp_src_endofpacket -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                           // limiter_001:rsp_src_valid -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                   // limiter_001:rsp_src_startofpacket -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [90:0] limiter_001_rsp_src_data;                                                                            // limiter_001:rsp_src_data -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [10:0] limiter_001_rsp_src_channel;                                                                         // limiter_001:rsp_src_channel -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                           // nios2_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         burst_adapter_source0_endofpacket;                                                                   // burst_adapter:source0_endofpacket -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                                         // burst_adapter:source0_valid -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                                 // burst_adapter:source0_startofpacket -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [63:0] burst_adapter_source0_data;                                                                          // burst_adapter:source0_data -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                                         // FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire  [10:0] burst_adapter_source0_channel;                                                                       // burst_adapter:source0_channel -> FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_001_source0_endofpacket;                                                               // burst_adapter_001:source0_endofpacket -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_001_source0_valid;                                                                     // burst_adapter_001:source0_valid -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_001_source0_startofpacket;                                                             // burst_adapter_001:source0_startofpacket -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [63:0] burst_adapter_001_source0_data;                                                                      // burst_adapter_001:source0_data -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_001_source0_ready;                                                                     // KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire  [10:0] burst_adapter_001_source0_channel;                                                                   // burst_adapter_001:source0_channel -> KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_002_source0_endofpacket;                                                               // burst_adapter_002:source0_endofpacket -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_002_source0_valid;                                                                     // burst_adapter_002:source0_valid -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_002_source0_startofpacket;                                                             // burst_adapter_002:source0_startofpacket -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [63:0] burst_adapter_002_source0_data;                                                                      // burst_adapter_002:source0_data -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_002_source0_ready;                                                                     // Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire  [10:0] burst_adapter_002_source0_channel;                                                                   // burst_adapter_002:source0_channel -> Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_003_source0_endofpacket;                                                               // burst_adapter_003:source0_endofpacket -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_003_source0_valid;                                                                     // burst_adapter_003:source0_valid -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_003_source0_startofpacket;                                                             // burst_adapter_003:source0_startofpacket -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [63:0] burst_adapter_003_source0_data;                                                                      // burst_adapter_003:source0_data -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_003_source0_ready;                                                                     // Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire  [10:0] burst_adapter_003_source0_channel;                                                                   // burst_adapter_003:source0_channel -> Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rst_controller_reset_out_reset;                                                                      // rst_controller:reset_out -> [FreqSynth_IP_0:reset_n, FreqSynth_IP_0_avalon_slave_0_translator:reset, FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, FreqSynth_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Hex_Driver_IP_0:reset_n, Hex_Driver_IP_0_avalon_slave_0_translator:reset, Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Hex_Driver_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Ir_Decode_IP_0:reset_n, Ir_Decode_IP_0_avalon_slave_0_translator:reset, Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Ir_Decode_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, KeyBoard_IP_0:reset_n, KeyBoard_IP_0_avalon_slave_0_translator:reset, KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, KeyBoard_IP_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, nios2:reset_n, nios2_data_master_translator:reset, nios2_data_master_translator_avalon_universal_master_0_agent:reset, nios2_instruction_master_translator:reset, nios2_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_jtag_debug_module_translator:reset, nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_led:reset_n, pio_led_s1_translator:reset, pio_led_s1_translator_avalon_universal_slave_0_agent:reset, pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ram:reset, ram_s1_translator:reset, ram_s1_translator_avalon_universal_slave_0_agent:reset, ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rom:reset, rom_s1_translator:reset, rom_s1_translator_avalon_universal_slave_0_agent:reset, rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset]
	wire         nios2_jtag_debug_module_reset_reset;                                                                 // nios2:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         cmd_xbar_demux_src0_endofpacket;                                                                     // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                           // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                   // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [90:0] cmd_xbar_demux_src0_data;                                                                            // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [10:0] cmd_xbar_demux_src0_channel;                                                                         // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                           // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                     // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                           // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                   // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [90:0] cmd_xbar_demux_src1_data;                                                                            // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [10:0] cmd_xbar_demux_src1_channel;                                                                         // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                           // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                     // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                           // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                   // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [90:0] cmd_xbar_demux_src2_data;                                                                            // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire  [10:0] cmd_xbar_demux_src2_channel;                                                                         // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                           // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                 // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                       // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                               // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [90:0] cmd_xbar_demux_001_src0_data;                                                                        // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [10:0] cmd_xbar_demux_001_src0_channel;                                                                     // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                       // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                 // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                       // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                               // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [90:0] cmd_xbar_demux_001_src1_data;                                                                        // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [10:0] cmd_xbar_demux_001_src1_channel;                                                                     // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                       // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                 // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                       // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                               // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [90:0] cmd_xbar_demux_001_src2_data;                                                                        // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire  [10:0] cmd_xbar_demux_001_src2_channel;                                                                     // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                       // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                 // cmd_xbar_demux_001:src3_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                       // cmd_xbar_demux_001:src3_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                               // cmd_xbar_demux_001:src3_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [90:0] cmd_xbar_demux_001_src3_data;                                                                        // cmd_xbar_demux_001:src3_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [10:0] cmd_xbar_demux_001_src3_channel;                                                                     // cmd_xbar_demux_001:src3_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                 // cmd_xbar_demux_001:src4_endofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                       // cmd_xbar_demux_001:src4_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                               // cmd_xbar_demux_001:src4_startofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [90:0] cmd_xbar_demux_001_src4_data;                                                                        // cmd_xbar_demux_001:src4_data -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [10:0] cmd_xbar_demux_001_src4_channel;                                                                     // cmd_xbar_demux_001:src4_channel -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                 // cmd_xbar_demux_001:src5_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                       // cmd_xbar_demux_001:src5_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                               // cmd_xbar_demux_001:src5_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [90:0] cmd_xbar_demux_001_src5_data;                                                                        // cmd_xbar_demux_001:src5_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [10:0] cmd_xbar_demux_001_src5_channel;                                                                     // cmd_xbar_demux_001:src5_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                 // cmd_xbar_demux_001:src6_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                       // cmd_xbar_demux_001:src6_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                               // cmd_xbar_demux_001:src6_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [90:0] cmd_xbar_demux_001_src6_data;                                                                        // cmd_xbar_demux_001:src6_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [10:0] cmd_xbar_demux_001_src6_channel;                                                                     // cmd_xbar_demux_001:src6_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                 // cmd_xbar_demux_001:src7_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                       // cmd_xbar_demux_001:src7_valid -> width_adapter:in_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                               // cmd_xbar_demux_001:src7_startofpacket -> width_adapter:in_startofpacket
	wire  [90:0] cmd_xbar_demux_001_src7_data;                                                                        // cmd_xbar_demux_001:src7_data -> width_adapter:in_data
	wire  [10:0] cmd_xbar_demux_001_src7_channel;                                                                     // cmd_xbar_demux_001:src7_channel -> width_adapter:in_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                 // cmd_xbar_demux_001:src8_endofpacket -> width_adapter_002:in_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                       // cmd_xbar_demux_001:src8_valid -> width_adapter_002:in_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                               // cmd_xbar_demux_001:src8_startofpacket -> width_adapter_002:in_startofpacket
	wire  [90:0] cmd_xbar_demux_001_src8_data;                                                                        // cmd_xbar_demux_001:src8_data -> width_adapter_002:in_data
	wire  [10:0] cmd_xbar_demux_001_src8_channel;                                                                     // cmd_xbar_demux_001:src8_channel -> width_adapter_002:in_channel
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                                 // cmd_xbar_demux_001:src9_endofpacket -> width_adapter_004:in_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                       // cmd_xbar_demux_001:src9_valid -> width_adapter_004:in_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                               // cmd_xbar_demux_001:src9_startofpacket -> width_adapter_004:in_startofpacket
	wire  [90:0] cmd_xbar_demux_001_src9_data;                                                                        // cmd_xbar_demux_001:src9_data -> width_adapter_004:in_data
	wire  [10:0] cmd_xbar_demux_001_src9_channel;                                                                     // cmd_xbar_demux_001:src9_channel -> width_adapter_004:in_channel
	wire         cmd_xbar_demux_001_src10_endofpacket;                                                                // cmd_xbar_demux_001:src10_endofpacket -> width_adapter_006:in_endofpacket
	wire         cmd_xbar_demux_001_src10_valid;                                                                      // cmd_xbar_demux_001:src10_valid -> width_adapter_006:in_valid
	wire         cmd_xbar_demux_001_src10_startofpacket;                                                              // cmd_xbar_demux_001:src10_startofpacket -> width_adapter_006:in_startofpacket
	wire  [90:0] cmd_xbar_demux_001_src10_data;                                                                       // cmd_xbar_demux_001:src10_data -> width_adapter_006:in_data
	wire  [10:0] cmd_xbar_demux_001_src10_channel;                                                                    // cmd_xbar_demux_001:src10_channel -> width_adapter_006:in_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                     // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                           // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                   // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [90:0] rsp_xbar_demux_src0_data;                                                                            // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [10:0] rsp_xbar_demux_src0_channel;                                                                         // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                           // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                     // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                           // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                   // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [90:0] rsp_xbar_demux_src1_data;                                                                            // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [10:0] rsp_xbar_demux_src1_channel;                                                                         // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                           // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                 // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                       // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                               // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [90:0] rsp_xbar_demux_001_src0_data;                                                                        // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [10:0] rsp_xbar_demux_001_src0_channel;                                                                     // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                       // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                 // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                       // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                               // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [90:0] rsp_xbar_demux_001_src1_data;                                                                        // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [10:0] rsp_xbar_demux_001_src1_channel;                                                                     // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                       // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                 // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                       // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                               // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [90:0] rsp_xbar_demux_002_src0_data;                                                                        // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [10:0] rsp_xbar_demux_002_src0_channel;                                                                     // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                       // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                 // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                       // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                               // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [90:0] rsp_xbar_demux_002_src1_data;                                                                        // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire  [10:0] rsp_xbar_demux_002_src1_channel;                                                                     // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                       // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                 // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                       // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                               // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [90:0] rsp_xbar_demux_003_src0_data;                                                                        // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire  [10:0] rsp_xbar_demux_003_src0_channel;                                                                     // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                       // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                 // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                       // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                               // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [90:0] rsp_xbar_demux_004_src0_data;                                                                        // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire  [10:0] rsp_xbar_demux_004_src0_channel;                                                                     // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                       // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                 // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                       // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                               // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [90:0] rsp_xbar_demux_005_src0_data;                                                                        // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire  [10:0] rsp_xbar_demux_005_src0_channel;                                                                     // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                       // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                 // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                       // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                               // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [90:0] rsp_xbar_demux_006_src0_data;                                                                        // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire  [10:0] rsp_xbar_demux_006_src0_channel;                                                                     // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                       // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                 // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                       // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                               // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [90:0] rsp_xbar_demux_007_src0_data;                                                                        // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire  [10:0] rsp_xbar_demux_007_src0_channel;                                                                     // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                       // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                 // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                       // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                               // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [90:0] rsp_xbar_demux_008_src0_data;                                                                        // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire  [10:0] rsp_xbar_demux_008_src0_channel;                                                                     // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                       // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                                 // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                       // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                               // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [90:0] rsp_xbar_demux_009_src0_data;                                                                        // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire  [10:0] rsp_xbar_demux_009_src0_channel;                                                                     // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                       // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                                 // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                       // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                               // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [90:0] rsp_xbar_demux_010_src0_data;                                                                        // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire  [10:0] rsp_xbar_demux_010_src0_channel;                                                                     // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                       // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                         // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                       // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [90:0] limiter_cmd_src_data;                                                                                // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire  [10:0] limiter_cmd_src_channel;                                                                             // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                               // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                        // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                              // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                      // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [90:0] rsp_xbar_mux_src_data;                                                                               // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire  [10:0] rsp_xbar_mux_src_channel;                                                                            // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                              // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                     // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                   // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [90:0] limiter_001_cmd_src_data;                                                                            // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire  [10:0] limiter_001_cmd_src_channel;                                                                         // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                           // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                    // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                          // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                  // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [90:0] rsp_xbar_mux_001_src_data;                                                                           // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire  [10:0] rsp_xbar_mux_001_src_channel;                                                                        // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                          // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                        // cmd_xbar_mux:src_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                              // cmd_xbar_mux:src_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                      // cmd_xbar_mux:src_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [90:0] cmd_xbar_mux_src_data;                                                                               // cmd_xbar_mux:src_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [10:0] cmd_xbar_mux_src_channel;                                                                            // cmd_xbar_mux:src_channel -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                              // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                           // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                 // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                         // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [90:0] id_router_src_data;                                                                                  // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [10:0] id_router_src_channel;                                                                               // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                 // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                    // cmd_xbar_mux_001:src_endofpacket -> rom_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                          // cmd_xbar_mux_001:src_valid -> rom_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                  // cmd_xbar_mux_001:src_startofpacket -> rom_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [90:0] cmd_xbar_mux_001_src_data;                                                                           // cmd_xbar_mux_001:src_data -> rom_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [10:0] cmd_xbar_mux_001_src_channel;                                                                        // cmd_xbar_mux_001:src_channel -> rom_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                          // rom_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                       // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                             // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                     // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [90:0] id_router_001_src_data;                                                                              // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [10:0] id_router_001_src_channel;                                                                           // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                             // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                    // cmd_xbar_mux_002:src_endofpacket -> ram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                          // cmd_xbar_mux_002:src_valid -> ram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                  // cmd_xbar_mux_002:src_startofpacket -> ram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [90:0] cmd_xbar_mux_002_src_data;                                                                           // cmd_xbar_mux_002:src_data -> ram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [10:0] cmd_xbar_mux_002_src_channel;                                                                        // cmd_xbar_mux_002:src_channel -> ram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                          // ram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                       // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                             // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                     // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [90:0] id_router_002_src_data;                                                                              // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [10:0] id_router_002_src_channel;                                                                           // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                             // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                                       // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                             // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                     // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [90:0] id_router_003_src_data;                                                                              // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [10:0] id_router_003_src_channel;                                                                           // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                             // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                       // pio_led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                       // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                             // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                     // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [90:0] id_router_004_src_data;                                                                              // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [10:0] id_router_004_src_channel;                                                                           // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                             // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                       // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                             // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                     // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [90:0] id_router_005_src_data;                                                                              // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [10:0] id_router_005_src_channel;                                                                           // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                             // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                                       // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                             // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                     // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [90:0] id_router_006_src_data;                                                                              // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [10:0] id_router_006_src_channel;                                                                           // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                             // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                                       // width_adapter:in_ready -> cmd_xbar_demux_001:src7_ready
	wire         width_adapter_src_endofpacket;                                                                       // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                             // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire         width_adapter_src_startofpacket;                                                                     // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [63:0] width_adapter_src_data;                                                                              // width_adapter:out_data -> burst_adapter:sink0_data
	wire         width_adapter_src_ready;                                                                             // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire  [10:0] width_adapter_src_channel;                                                                           // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire         id_router_007_src_endofpacket;                                                                       // id_router_007:src_endofpacket -> width_adapter_001:in_endofpacket
	wire         id_router_007_src_valid;                                                                             // id_router_007:src_valid -> width_adapter_001:in_valid
	wire         id_router_007_src_startofpacket;                                                                     // id_router_007:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [63:0] id_router_007_src_data;                                                                              // id_router_007:src_data -> width_adapter_001:in_data
	wire  [10:0] id_router_007_src_channel;                                                                           // id_router_007:src_channel -> width_adapter_001:in_channel
	wire         id_router_007_src_ready;                                                                             // width_adapter_001:in_ready -> id_router_007:src_ready
	wire         width_adapter_001_src_endofpacket;                                                                   // width_adapter_001:out_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         width_adapter_001_src_valid;                                                                         // width_adapter_001:out_valid -> rsp_xbar_demux_007:sink_valid
	wire         width_adapter_001_src_startofpacket;                                                                 // width_adapter_001:out_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [90:0] width_adapter_001_src_data;                                                                          // width_adapter_001:out_data -> rsp_xbar_demux_007:sink_data
	wire         width_adapter_001_src_ready;                                                                         // rsp_xbar_demux_007:sink_ready -> width_adapter_001:out_ready
	wire  [10:0] width_adapter_001_src_channel;                                                                       // width_adapter_001:out_channel -> rsp_xbar_demux_007:sink_channel
	wire         cmd_xbar_demux_001_src8_ready;                                                                       // width_adapter_002:in_ready -> cmd_xbar_demux_001:src8_ready
	wire         width_adapter_002_src_endofpacket;                                                                   // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire         width_adapter_002_src_valid;                                                                         // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire         width_adapter_002_src_startofpacket;                                                                 // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [63:0] width_adapter_002_src_data;                                                                          // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire         width_adapter_002_src_ready;                                                                         // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire  [10:0] width_adapter_002_src_channel;                                                                       // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire         id_router_008_src_endofpacket;                                                                       // id_router_008:src_endofpacket -> width_adapter_003:in_endofpacket
	wire         id_router_008_src_valid;                                                                             // id_router_008:src_valid -> width_adapter_003:in_valid
	wire         id_router_008_src_startofpacket;                                                                     // id_router_008:src_startofpacket -> width_adapter_003:in_startofpacket
	wire  [63:0] id_router_008_src_data;                                                                              // id_router_008:src_data -> width_adapter_003:in_data
	wire  [10:0] id_router_008_src_channel;                                                                           // id_router_008:src_channel -> width_adapter_003:in_channel
	wire         id_router_008_src_ready;                                                                             // width_adapter_003:in_ready -> id_router_008:src_ready
	wire         width_adapter_003_src_endofpacket;                                                                   // width_adapter_003:out_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         width_adapter_003_src_valid;                                                                         // width_adapter_003:out_valid -> rsp_xbar_demux_008:sink_valid
	wire         width_adapter_003_src_startofpacket;                                                                 // width_adapter_003:out_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [90:0] width_adapter_003_src_data;                                                                          // width_adapter_003:out_data -> rsp_xbar_demux_008:sink_data
	wire         width_adapter_003_src_ready;                                                                         // rsp_xbar_demux_008:sink_ready -> width_adapter_003:out_ready
	wire  [10:0] width_adapter_003_src_channel;                                                                       // width_adapter_003:out_channel -> rsp_xbar_demux_008:sink_channel
	wire         cmd_xbar_demux_001_src9_ready;                                                                       // width_adapter_004:in_ready -> cmd_xbar_demux_001:src9_ready
	wire         width_adapter_004_src_endofpacket;                                                                   // width_adapter_004:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire         width_adapter_004_src_valid;                                                                         // width_adapter_004:out_valid -> burst_adapter_002:sink0_valid
	wire         width_adapter_004_src_startofpacket;                                                                 // width_adapter_004:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire  [63:0] width_adapter_004_src_data;                                                                          // width_adapter_004:out_data -> burst_adapter_002:sink0_data
	wire         width_adapter_004_src_ready;                                                                         // burst_adapter_002:sink0_ready -> width_adapter_004:out_ready
	wire  [10:0] width_adapter_004_src_channel;                                                                       // width_adapter_004:out_channel -> burst_adapter_002:sink0_channel
	wire         id_router_009_src_endofpacket;                                                                       // id_router_009:src_endofpacket -> width_adapter_005:in_endofpacket
	wire         id_router_009_src_valid;                                                                             // id_router_009:src_valid -> width_adapter_005:in_valid
	wire         id_router_009_src_startofpacket;                                                                     // id_router_009:src_startofpacket -> width_adapter_005:in_startofpacket
	wire  [63:0] id_router_009_src_data;                                                                              // id_router_009:src_data -> width_adapter_005:in_data
	wire  [10:0] id_router_009_src_channel;                                                                           // id_router_009:src_channel -> width_adapter_005:in_channel
	wire         id_router_009_src_ready;                                                                             // width_adapter_005:in_ready -> id_router_009:src_ready
	wire         width_adapter_005_src_endofpacket;                                                                   // width_adapter_005:out_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         width_adapter_005_src_valid;                                                                         // width_adapter_005:out_valid -> rsp_xbar_demux_009:sink_valid
	wire         width_adapter_005_src_startofpacket;                                                                 // width_adapter_005:out_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [90:0] width_adapter_005_src_data;                                                                          // width_adapter_005:out_data -> rsp_xbar_demux_009:sink_data
	wire         width_adapter_005_src_ready;                                                                         // rsp_xbar_demux_009:sink_ready -> width_adapter_005:out_ready
	wire  [10:0] width_adapter_005_src_channel;                                                                       // width_adapter_005:out_channel -> rsp_xbar_demux_009:sink_channel
	wire         cmd_xbar_demux_001_src10_ready;                                                                      // width_adapter_006:in_ready -> cmd_xbar_demux_001:src10_ready
	wire         width_adapter_006_src_endofpacket;                                                                   // width_adapter_006:out_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire         width_adapter_006_src_valid;                                                                         // width_adapter_006:out_valid -> burst_adapter_003:sink0_valid
	wire         width_adapter_006_src_startofpacket;                                                                 // width_adapter_006:out_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire  [63:0] width_adapter_006_src_data;                                                                          // width_adapter_006:out_data -> burst_adapter_003:sink0_data
	wire         width_adapter_006_src_ready;                                                                         // burst_adapter_003:sink0_ready -> width_adapter_006:out_ready
	wire  [10:0] width_adapter_006_src_channel;                                                                       // width_adapter_006:out_channel -> burst_adapter_003:sink0_channel
	wire         id_router_010_src_endofpacket;                                                                       // id_router_010:src_endofpacket -> width_adapter_007:in_endofpacket
	wire         id_router_010_src_valid;                                                                             // id_router_010:src_valid -> width_adapter_007:in_valid
	wire         id_router_010_src_startofpacket;                                                                     // id_router_010:src_startofpacket -> width_adapter_007:in_startofpacket
	wire  [63:0] id_router_010_src_data;                                                                              // id_router_010:src_data -> width_adapter_007:in_data
	wire  [10:0] id_router_010_src_channel;                                                                           // id_router_010:src_channel -> width_adapter_007:in_channel
	wire         id_router_010_src_ready;                                                                             // width_adapter_007:in_ready -> id_router_010:src_ready
	wire         width_adapter_007_src_endofpacket;                                                                   // width_adapter_007:out_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         width_adapter_007_src_valid;                                                                         // width_adapter_007:out_valid -> rsp_xbar_demux_010:sink_valid
	wire         width_adapter_007_src_startofpacket;                                                                 // width_adapter_007:out_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [90:0] width_adapter_007_src_data;                                                                          // width_adapter_007:out_data -> rsp_xbar_demux_010:sink_data
	wire         width_adapter_007_src_ready;                                                                         // rsp_xbar_demux_010:sink_ready -> width_adapter_007:out_ready
	wire  [10:0] width_adapter_007_src_channel;                                                                       // width_adapter_007:out_channel -> rsp_xbar_demux_010:sink_channel
	wire  [10:0] limiter_cmd_valid_data;                                                                              // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire  [10:0] limiter_001_cmd_valid_data;                                                                          // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                            // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                            // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_d_irq_irq;                                                                                     // irq_mapper:sender_irq -> nios2:d_irq

	mysystem_nios2 nios2 (
		.clk                                   (clk_clk),                                                            //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                    //                   reset_n.reset_n
		.d_address                             (nios2_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_data_master_writedata),                                        //                          .writedata
		.d_readdatavalid                       (nios2_data_master_readdatavalid),                                    //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (nios2_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (nios2_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	mysystem_rom rom (
		.clk         (clk_clk),                                           //   clk1.clk
		.address     (rom_s1_translator_avalon_anti_slave_0_address),     //     s1.address
		.debugaccess (rom_s1_translator_avalon_anti_slave_0_debugaccess), //       .debugaccess
		.clken       (rom_s1_translator_avalon_anti_slave_0_clken),       //       .clken
		.chipselect  (rom_s1_translator_avalon_anti_slave_0_chipselect),  //       .chipselect
		.write       (rom_s1_translator_avalon_anti_slave_0_write),       //       .write
		.readdata    (rom_s1_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.writedata   (rom_s1_translator_avalon_anti_slave_0_writedata),   //       .writedata
		.byteenable  (rom_s1_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset)                     // reset1.reset
	);

	mysystem_ram ram (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (ram_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (ram_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (ram_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (ram_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (ram_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (ram_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ram_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                    // reset1.reset
	);

	mysystem_sysid sysid (
		.clock    (clk_clk),                                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                             //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	mysystem_pio_led pio_led (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (pio_led_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_led_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_led_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_led_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_led_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_export)                                            // external_connection.export
	);

	mysystem_timer_0 timer_0 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                              //   irq.irq
	);

	mysystem_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                  //               irq.irq
	);

	avalon_FreqSynth freqsynth_ip_0 (
		.clk        (clk_clk),                                                                 //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                                         //          reset.reset_n
		.address    (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    // avalon_slave_0.address
		.writedata  (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.write      (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.read       (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.chipselect (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.readdata   (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.vib        (vib_export_export)                                                        //    conduit_end.export
	);

	avalon_KeyBoard keyboard_ip_0 (
		.clk             (clk_clk),                                                                //          clock.clk
		.reset_n         (~rst_controller_reset_out_reset),                                        //          reset.reset_n
		.address         (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    // avalon_slave_0.address
		.read            (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.chipselect      (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.readdata        (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata       (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.write           (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.Key_Board_Row_i (keyboard_export_Row_i),                                                  //    conduit_end.export
		.Key_Board_Col_o (keyboard_export_Col_o)                                                   //               .export
	);

	avalon_ir_decode ir_decode_ip_0 (
		.clk        (clk_clk),                                                                 //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                                         //          reset.reset_n
		.address    (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    // avalon_slave_0.address
		.writedata  (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.write      (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.read       (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.chipselect (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.readdata   (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.iIR        (ir_decode_export_iIR),                                                    //    conduit_end.export
		.Get_Flag_o (ir_decode_export_Get_Flag_o)                                              //               .export
	);

	avalon_hex_top hex_driver_ip_0 (
		.clk        (clk_clk),                                                                  //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                                          //          reset.reset_n
		.address    (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    // avalon_slave_0.address
		.writedata  (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.write      (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.read       (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.chipselect (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.readdata   (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.SH_CP      (hex_driver_export_SH_CP),                                                  //    conduit_end.export
		.ST_CP      (hex_driver_export_ST_CP),                                                  //               .export
		.DS         (hex_driver_export_DS)                                                      //               .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_instruction_master_translator (
		.clk                      (clk_clk),                                                                     //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (nios2_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_byteenable            (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_write                 (1'b0),                                                                        //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.av_debugaccess           (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_data_master_translator (
		.clk                      (clk_clk),                                                              //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address              (nios2_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_data_master_read),                                               //                          .read
		.av_readdata              (nios2_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (nios2_data_master_write),                                              //                          .write
		.av_writedata             (nios2_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                 //               (terminated)
		.av_begintransfer         (1'b0),                                                                 //               (terminated)
		.av_chipselect            (1'b0),                                                                 //               (terminated)
		.av_lock                  (1'b0),                                                                 //               (terminated)
		.uav_clken                (),                                                                     //               (terminated)
		.av_clken                 (1'b1),                                                                 //               (terminated)
		.uav_response             (2'b00),                                                                //               (terminated)
		.av_response              (),                                                                     //               (terminated)
		.uav_writeresponserequest (),                                                                     //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                 //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                 //               (terminated)
		.av_writeresponsevalid    ()                                                                      //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_chipselect            (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rom_s1_translator (
		.clk                      (clk_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address              (rom_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (rom_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (rom_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (rom_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (rom_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (rom_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (rom_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (rom_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (rom_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (rom_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (rom_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (rom_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (rom_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (rom_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (rom_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (rom_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (rom_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (rom_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_debugaccess           (rom_s1_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ram_s1_translator (
		.clk                      (clk_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address              (ram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (ram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (ram_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_led_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_led_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_led_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_led_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_led_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_led_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) freqsynth_ip_0_avalon_slave_0_translator (
		.clk                      (clk_clk),                                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (freqsynth_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) keyboard_ip_0_avalon_slave_0_translator (
		.clk                      (clk_clk),                                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address              (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (keyboard_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                                        //              (terminated)
		.av_burstcount            (),                                                                                        //              (terminated)
		.av_byteenable            (),                                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                                        //              (terminated)
		.av_lock                  (),                                                                                        //              (terminated)
		.av_clken                 (),                                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                                    //              (terminated)
		.av_debugaccess           (),                                                                                        //              (terminated)
		.av_outputenable          (),                                                                                        //              (terminated)
		.uav_response             (),                                                                                        //              (terminated)
		.av_response              (2'b00),                                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ir_decode_ip_0_avalon_slave_0_translator (
		.clk                      (clk_clk),                                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ir_decode_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex_driver_ip_0_avalon_slave_0_translator (
		.clk                      (clk_clk),                                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex_driver_ip_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_byteenable            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_debugaccess           (),                                                                                          //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_THREAD_ID_H           (81),
		.PKT_THREAD_ID_L           (81),
		.PKT_CACHE_H               (88),
		.PKT_CACHE_L               (85),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                              //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (nios2_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                                //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                                 //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                              //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                        //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                          //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                                //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_THREAD_ID_H           (81),
		.PKT_THREAD_ID_L           (81),
		.PKT_CACHE_H               (88),
		.PKT_CACHE_L               (85),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                       //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address              (nios2_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                     //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                      //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                                   //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                             //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                               //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                     //          .ready
		.av_response             (),                                                                              // (terminated)
		.av_writeresponserequest (1'b0),                                                                          // (terminated)
		.av_writeresponsevalid   ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                     //                .channel
		.rf_sink_ready           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) rom_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (rom_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rom_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rom_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rom_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rom_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rom_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rom_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rom_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rom_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rom_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rom_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rom_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rom_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rom_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rom_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rom_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                //                .channel
		.rf_sink_ready           (rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rom_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rom_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rom_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rom_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rom_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (rom_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rom_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rom_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rom_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rom_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (ram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                //                .channel
		.rf_sink_ready           (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_led_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                 //                .channel
		.rf_sink_ready           (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                 //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (44),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (24),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (25),
		.PKT_TRANS_POSTED          (26),
		.PKT_TRANS_WRITE           (27),
		.PKT_TRANS_READ            (28),
		.PKT_TRANS_LOCK            (29),
		.PKT_SRC_ID_H              (49),
		.PKT_SRC_ID_L              (46),
		.PKT_DEST_ID_H             (53),
		.PKT_DEST_ID_L             (50),
		.PKT_BURSTWRAP_H           (36),
		.PKT_BURSTWRAP_L           (34),
		.PKT_BYTE_CNT_H            (33),
		.PKT_BYTE_CNT_L            (31),
		.PKT_PROTECTION_H          (57),
		.PKT_PROTECTION_L          (55),
		.PKT_RESPONSE_STATUS_H     (63),
		.PKT_RESPONSE_STATUS_L     (62),
		.PKT_BURST_SIZE_H          (39),
		.PKT_BURST_SIZE_L          (37),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (64),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                        //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                        //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                         //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                                      //                .channel
		.rf_sink_ready           (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (65),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (44),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (24),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (25),
		.PKT_TRANS_POSTED          (26),
		.PKT_TRANS_WRITE           (27),
		.PKT_TRANS_READ            (28),
		.PKT_TRANS_LOCK            (29),
		.PKT_SRC_ID_H              (49),
		.PKT_SRC_ID_L              (46),
		.PKT_DEST_ID_H             (53),
		.PKT_DEST_ID_L             (50),
		.PKT_BURSTWRAP_H           (36),
		.PKT_BURSTWRAP_L           (34),
		.PKT_BYTE_CNT_H            (33),
		.PKT_BYTE_CNT_L            (31),
		.PKT_PROTECTION_H          (57),
		.PKT_PROTECTION_L          (55),
		.PKT_RESPONSE_STATUS_H     (63),
		.PKT_RESPONSE_STATUS_L     (62),
		.PKT_BURST_SIZE_H          (39),
		.PKT_BURST_SIZE_L          (37),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (64),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                                   //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                                   //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                                    //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                             //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                                 //                .channel
		.rf_sink_ready           (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (65),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (44),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (24),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (25),
		.PKT_TRANS_POSTED          (26),
		.PKT_TRANS_WRITE           (27),
		.PKT_TRANS_READ            (28),
		.PKT_TRANS_LOCK            (29),
		.PKT_SRC_ID_H              (49),
		.PKT_SRC_ID_L              (46),
		.PKT_DEST_ID_H             (53),
		.PKT_DEST_ID_L             (50),
		.PKT_BURSTWRAP_H           (36),
		.PKT_BURSTWRAP_L           (34),
		.PKT_BYTE_CNT_H            (33),
		.PKT_BYTE_CNT_L            (31),
		.PKT_PROTECTION_H          (57),
		.PKT_PROTECTION_L          (55),
		.PKT_RESPONSE_STATUS_H     (63),
		.PKT_RESPONSE_STATUS_L     (62),
		.PKT_BURST_SIZE_H          (39),
		.PKT_BURST_SIZE_L          (37),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (64),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                                    //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                                    //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                                     //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                              //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                                  //                .channel
		.rf_sink_ready           (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (65),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (44),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (24),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (25),
		.PKT_TRANS_POSTED          (26),
		.PKT_TRANS_WRITE           (27),
		.PKT_TRANS_READ            (28),
		.PKT_TRANS_LOCK            (29),
		.PKT_SRC_ID_H              (49),
		.PKT_SRC_ID_L              (46),
		.PKT_DEST_ID_H             (53),
		.PKT_DEST_ID_L             (50),
		.PKT_BURSTWRAP_H           (36),
		.PKT_BURSTWRAP_L           (34),
		.PKT_BYTE_CNT_H            (33),
		.PKT_BYTE_CNT_L            (31),
		.PKT_PROTECTION_H          (57),
		.PKT_PROTECTION_L          (55),
		.PKT_RESPONSE_STATUS_H     (63),
		.PKT_RESPONSE_STATUS_L     (62),
		.PKT_BURST_SIZE_H          (39),
		.PKT_BURST_SIZE_L          (37),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (64),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                                     //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                                     //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                                      //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                               //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                                   //                .channel
		.rf_sink_ready           (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (65),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	mysystem_addr_router addr_router (
		.sink_ready         (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	mysystem_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                     //          .valid
		.src_data           (addr_router_001_src_data),                                                      //          .data
		.src_channel        (addr_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                //          .endofpacket
	);

	mysystem_id_router id_router (
		.sink_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                //       src.ready
		.src_valid          (id_router_src_valid),                                                                //          .valid
		.src_data           (id_router_src_data),                                                                 //          .data
		.src_channel        (id_router_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                           //          .endofpacket
	);

	mysystem_id_router id_router_001 (
		.sink_ready         (rom_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rom_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rom_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rom_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rom_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                           //       src.ready
		.src_valid          (id_router_001_src_valid),                                           //          .valid
		.src_data           (id_router_001_src_data),                                            //          .data
		.src_channel        (id_router_001_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                      //          .endofpacket
	);

	mysystem_id_router id_router_002 (
		.sink_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                           //       src.ready
		.src_valid          (id_router_002_src_valid),                                           //          .valid
		.src_data           (id_router_002_src_data),                                            //          .data
		.src_channel        (id_router_002_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                      //          .endofpacket
	);

	mysystem_id_router_003 id_router_003 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                        //       src.ready
		.src_valid          (id_router_003_src_valid),                                                        //          .valid
		.src_data           (id_router_003_src_data),                                                         //          .data
		.src_channel        (id_router_003_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                   //          .endofpacket
	);

	mysystem_id_router_003 id_router_004 (
		.sink_ready         (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                               //       src.ready
		.src_valid          (id_router_004_src_valid),                                               //          .valid
		.src_data           (id_router_004_src_data),                                                //          .data
		.src_channel        (id_router_004_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                          //          .endofpacket
	);

	mysystem_id_router_003 id_router_005 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                               //       src.ready
		.src_valid          (id_router_005_src_valid),                                               //          .valid
		.src_data           (id_router_005_src_data),                                                //          .data
		.src_channel        (id_router_005_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                          //          .endofpacket
	);

	mysystem_id_router_003 id_router_006 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                  //          .valid
		.src_data           (id_router_006_src_data),                                                                   //          .data
		.src_channel        (id_router_006_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                             //          .endofpacket
	);

	mysystem_id_router_007 id_router_007 (
		.sink_ready         (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (freqsynth_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_007_src_valid),                                                                  //          .valid
		.src_data           (id_router_007_src_data),                                                                   //          .data
		.src_channel        (id_router_007_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                             //          .endofpacket
	);

	mysystem_id_router_007 id_router_008 (
		.sink_ready         (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (keyboard_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                 //          .valid
		.src_data           (id_router_008_src_data),                                                                  //          .data
		.src_channel        (id_router_008_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                            //          .endofpacket
	);

	mysystem_id_router_007 id_router_009 (
		.sink_ready         (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ir_decode_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_009_src_valid),                                                                  //          .valid
		.src_data           (id_router_009_src_data),                                                                   //          .data
		.src_channel        (id_router_009_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                             //          .endofpacket
	);

	mysystem_id_router_007 id_router_010 (
		.sink_ready         (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex_driver_ip_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_010_src_valid),                                                                   //          .valid
		.src_data           (id_router_010_src_data),                                                                    //          .data
		.src_channel        (id_router_010_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                              //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (11),
		.VALID_WIDTH               (11),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.MAX_OUTSTANDING_RESPONSES (3),
		.PIPELINED                 (0),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (11),
		.VALID_WIDTH               (11),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (24),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (44),
		.PKT_BYTE_CNT_H            (33),
		.PKT_BYTE_CNT_L            (31),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (39),
		.PKT_BURST_SIZE_L          (37),
		.PKT_BURST_TYPE_H          (41),
		.PKT_BURST_TYPE_L          (40),
		.PKT_BURSTWRAP_H           (36),
		.PKT_BURSTWRAP_L           (34),
		.PKT_TRANS_COMPRESSED_READ (25),
		.PKT_TRANS_WRITE           (27),
		.PKT_TRANS_READ            (28),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (64),
		.ST_CHANNEL_W              (11),
		.OUT_BYTE_CNT_H            (31),
		.OUT_BURSTWRAP_H           (36),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter (
		.clk                   (clk_clk),                             //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (24),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (44),
		.PKT_BYTE_CNT_H            (33),
		.PKT_BYTE_CNT_L            (31),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (39),
		.PKT_BURST_SIZE_L          (37),
		.PKT_BURST_TYPE_H          (41),
		.PKT_BURST_TYPE_L          (40),
		.PKT_BURSTWRAP_H           (36),
		.PKT_BURSTWRAP_L           (34),
		.PKT_TRANS_COMPRESSED_READ (25),
		.PKT_TRANS_WRITE           (27),
		.PKT_TRANS_READ            (28),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (64),
		.ST_CHANNEL_W              (11),
		.OUT_BYTE_CNT_H            (31),
		.OUT_BURSTWRAP_H           (36),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_001 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (24),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (44),
		.PKT_BYTE_CNT_H            (33),
		.PKT_BYTE_CNT_L            (31),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (39),
		.PKT_BURST_SIZE_L          (37),
		.PKT_BURST_TYPE_H          (41),
		.PKT_BURST_TYPE_L          (40),
		.PKT_BURSTWRAP_H           (36),
		.PKT_BURSTWRAP_L           (34),
		.PKT_TRANS_COMPRESSED_READ (25),
		.PKT_TRANS_WRITE           (27),
		.PKT_TRANS_READ            (28),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (64),
		.ST_CHANNEL_W              (11),
		.OUT_BYTE_CNT_H            (31),
		.OUT_BURSTWRAP_H           (36),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_002 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (24),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (44),
		.PKT_BYTE_CNT_H            (33),
		.PKT_BYTE_CNT_L            (31),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (39),
		.PKT_BURST_SIZE_L          (37),
		.PKT_BURST_TYPE_H          (41),
		.PKT_BURST_TYPE_L          (40),
		.PKT_BURSTWRAP_H           (36),
		.PKT_BURSTWRAP_L           (34),
		.PKT_TRANS_COMPRESSED_READ (25),
		.PKT_TRANS_WRITE           (27),
		.PKT_TRANS_READ            (28),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (64),
		.ST_CHANNEL_W              (11),
		.OUT_BYTE_CNT_H            (31),
		.OUT_BURSTWRAP_H           (36),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_003 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_006_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_006_src_data),              //          .data
		.sink0_channel         (width_adapter_006_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_006_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_006_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_006_src_ready),             //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	mysystem_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //           .endofpacket
	);

	mysystem_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk_clk),                                //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket)    //           .endofpacket
	);

	mysystem_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	mysystem_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	mysystem_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_demux_003 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_demux_003 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_demux_003 rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_demux_003 rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_005_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_005_src_channel),         //          .channel
		.sink_data          (width_adapter_005_src_data),            //          .data
		.sink_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_005_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_demux_003 rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_007_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_007_src_channel),         //          .channel
		.sink_data          (width_adapter_007_src_data),            //          .data
		.sink_startofpacket (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_007_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	mysystem_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (51),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (60),
		.IN_PKT_BYTE_CNT_L             (58),
		.IN_PKT_TRANS_COMPRESSED_READ  (52),
		.IN_PKT_BURSTWRAP_H            (63),
		.IN_PKT_BURSTWRAP_L            (61),
		.IN_PKT_BURST_SIZE_H           (66),
		.IN_PKT_BURST_SIZE_L           (64),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (57),
		.IN_PKT_BURST_TYPE_H           (68),
		.IN_PKT_BURST_TYPE_L           (67),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (24),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (33),
		.OUT_PKT_BYTE_CNT_L            (31),
		.OUT_PKT_TRANS_COMPRESSED_READ (25),
		.OUT_PKT_BURST_SIZE_H          (39),
		.OUT_PKT_BURST_SIZE_L          (37),
		.OUT_PKT_RESPONSE_STATUS_H     (63),
		.OUT_PKT_RESPONSE_STATUS_L     (62),
		.OUT_PKT_TRANS_EXCLUSIVE       (30),
		.OUT_PKT_BURST_TYPE_H          (41),
		.OUT_PKT_BURST_TYPE_L          (40),
		.OUT_ST_DATA_W                 (64),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src7_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src7_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src7_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src7_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src7_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),         //       src.endofpacket
		.out_data             (width_adapter_src_data),                //          .data
		.out_channel          (width_adapter_src_channel),             //          .channel
		.out_valid            (width_adapter_src_valid),               //          .valid
		.out_ready            (width_adapter_src_ready),               //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),       //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (24),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (33),
		.IN_PKT_BYTE_CNT_L             (31),
		.IN_PKT_TRANS_COMPRESSED_READ  (25),
		.IN_PKT_BURSTWRAP_H            (36),
		.IN_PKT_BURSTWRAP_L            (34),
		.IN_PKT_BURST_SIZE_H           (39),
		.IN_PKT_BURST_SIZE_L           (37),
		.IN_PKT_RESPONSE_STATUS_H      (63),
		.IN_PKT_RESPONSE_STATUS_L      (62),
		.IN_PKT_TRANS_EXCLUSIVE        (30),
		.IN_PKT_BURST_TYPE_H           (41),
		.IN_PKT_BURST_TYPE_L           (40),
		.IN_ST_DATA_W                  (64),
		.OUT_PKT_ADDR_H                (51),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (60),
		.OUT_PKT_BYTE_CNT_L            (58),
		.OUT_PKT_TRANS_COMPRESSED_READ (52),
		.OUT_PKT_BURST_SIZE_H          (66),
		.OUT_PKT_BURST_SIZE_L          (64),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (57),
		.OUT_PKT_BURST_TYPE_H          (68),
		.OUT_PKT_BURST_TYPE_L          (67),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_007_src_valid),             //      sink.valid
		.in_channel           (id_router_007_src_channel),           //          .channel
		.in_startofpacket     (id_router_007_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_007_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_007_src_ready),             //          .ready
		.in_data              (id_router_007_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (51),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (60),
		.IN_PKT_BYTE_CNT_L             (58),
		.IN_PKT_TRANS_COMPRESSED_READ  (52),
		.IN_PKT_BURSTWRAP_H            (63),
		.IN_PKT_BURSTWRAP_L            (61),
		.IN_PKT_BURST_SIZE_H           (66),
		.IN_PKT_BURST_SIZE_L           (64),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (57),
		.IN_PKT_BURST_TYPE_H           (68),
		.IN_PKT_BURST_TYPE_L           (67),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (24),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (33),
		.OUT_PKT_BYTE_CNT_L            (31),
		.OUT_PKT_TRANS_COMPRESSED_READ (25),
		.OUT_PKT_BURST_SIZE_H          (39),
		.OUT_PKT_BURST_SIZE_L          (37),
		.OUT_PKT_RESPONSE_STATUS_H     (63),
		.OUT_PKT_RESPONSE_STATUS_L     (62),
		.OUT_PKT_TRANS_EXCLUSIVE       (30),
		.OUT_PKT_BURST_TYPE_H          (41),
		.OUT_PKT_BURST_TYPE_L          (40),
		.OUT_ST_DATA_W                 (64),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src8_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src8_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src8_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src8_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src8_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_002_src_data),            //          .data
		.out_channel          (width_adapter_002_src_channel),         //          .channel
		.out_valid            (width_adapter_002_src_valid),           //          .valid
		.out_ready            (width_adapter_002_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (24),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (33),
		.IN_PKT_BYTE_CNT_L             (31),
		.IN_PKT_TRANS_COMPRESSED_READ  (25),
		.IN_PKT_BURSTWRAP_H            (36),
		.IN_PKT_BURSTWRAP_L            (34),
		.IN_PKT_BURST_SIZE_H           (39),
		.IN_PKT_BURST_SIZE_L           (37),
		.IN_PKT_RESPONSE_STATUS_H      (63),
		.IN_PKT_RESPONSE_STATUS_L      (62),
		.IN_PKT_TRANS_EXCLUSIVE        (30),
		.IN_PKT_BURST_TYPE_H           (41),
		.IN_PKT_BURST_TYPE_L           (40),
		.IN_ST_DATA_W                  (64),
		.OUT_PKT_ADDR_H                (51),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (60),
		.OUT_PKT_BYTE_CNT_L            (58),
		.OUT_PKT_TRANS_COMPRESSED_READ (52),
		.OUT_PKT_BURST_SIZE_H          (66),
		.OUT_PKT_BURST_SIZE_L          (64),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (57),
		.OUT_PKT_BURST_TYPE_H          (68),
		.OUT_PKT_BURST_TYPE_L          (67),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_003 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_008_src_valid),             //      sink.valid
		.in_channel           (id_router_008_src_channel),           //          .channel
		.in_startofpacket     (id_router_008_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_008_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_008_src_ready),             //          .ready
		.in_data              (id_router_008_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (51),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (60),
		.IN_PKT_BYTE_CNT_L             (58),
		.IN_PKT_TRANS_COMPRESSED_READ  (52),
		.IN_PKT_BURSTWRAP_H            (63),
		.IN_PKT_BURSTWRAP_L            (61),
		.IN_PKT_BURST_SIZE_H           (66),
		.IN_PKT_BURST_SIZE_L           (64),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (57),
		.IN_PKT_BURST_TYPE_H           (68),
		.IN_PKT_BURST_TYPE_L           (67),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (24),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (33),
		.OUT_PKT_BYTE_CNT_L            (31),
		.OUT_PKT_TRANS_COMPRESSED_READ (25),
		.OUT_PKT_BURST_SIZE_H          (39),
		.OUT_PKT_BURST_SIZE_L          (37),
		.OUT_PKT_RESPONSE_STATUS_H     (63),
		.OUT_PKT_RESPONSE_STATUS_L     (62),
		.OUT_PKT_TRANS_EXCLUSIVE       (30),
		.OUT_PKT_BURST_TYPE_H          (41),
		.OUT_PKT_BURST_TYPE_L          (40),
		.OUT_ST_DATA_W                 (64),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_004 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src9_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src9_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src9_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src9_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src9_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_004_src_data),            //          .data
		.out_channel          (width_adapter_004_src_channel),         //          .channel
		.out_valid            (width_adapter_004_src_valid),           //          .valid
		.out_ready            (width_adapter_004_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (24),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (33),
		.IN_PKT_BYTE_CNT_L             (31),
		.IN_PKT_TRANS_COMPRESSED_READ  (25),
		.IN_PKT_BURSTWRAP_H            (36),
		.IN_PKT_BURSTWRAP_L            (34),
		.IN_PKT_BURST_SIZE_H           (39),
		.IN_PKT_BURST_SIZE_L           (37),
		.IN_PKT_RESPONSE_STATUS_H      (63),
		.IN_PKT_RESPONSE_STATUS_L      (62),
		.IN_PKT_TRANS_EXCLUSIVE        (30),
		.IN_PKT_BURST_TYPE_H           (41),
		.IN_PKT_BURST_TYPE_L           (40),
		.IN_ST_DATA_W                  (64),
		.OUT_PKT_ADDR_H                (51),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (60),
		.OUT_PKT_BYTE_CNT_L            (58),
		.OUT_PKT_TRANS_COMPRESSED_READ (52),
		.OUT_PKT_BURST_SIZE_H          (66),
		.OUT_PKT_BURST_SIZE_L          (64),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (57),
		.OUT_PKT_BURST_TYPE_H          (68),
		.OUT_PKT_BURST_TYPE_L          (67),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_005 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_009_src_valid),             //      sink.valid
		.in_channel           (id_router_009_src_channel),           //          .channel
		.in_startofpacket     (id_router_009_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_009_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_009_src_ready),             //          .ready
		.in_data              (id_router_009_src_data),              //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_005_src_data),          //          .data
		.out_channel          (width_adapter_005_src_channel),       //          .channel
		.out_valid            (width_adapter_005_src_valid),         //          .valid
		.out_ready            (width_adapter_005_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (51),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (60),
		.IN_PKT_BYTE_CNT_L             (58),
		.IN_PKT_TRANS_COMPRESSED_READ  (52),
		.IN_PKT_BURSTWRAP_H            (63),
		.IN_PKT_BURSTWRAP_L            (61),
		.IN_PKT_BURST_SIZE_H           (66),
		.IN_PKT_BURST_SIZE_L           (64),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (57),
		.IN_PKT_BURST_TYPE_H           (68),
		.IN_PKT_BURST_TYPE_L           (67),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (24),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (33),
		.OUT_PKT_BYTE_CNT_L            (31),
		.OUT_PKT_TRANS_COMPRESSED_READ (25),
		.OUT_PKT_BURST_SIZE_H          (39),
		.OUT_PKT_BURST_SIZE_L          (37),
		.OUT_PKT_RESPONSE_STATUS_H     (63),
		.OUT_PKT_RESPONSE_STATUS_L     (62),
		.OUT_PKT_TRANS_EXCLUSIVE       (30),
		.OUT_PKT_BURST_TYPE_H          (41),
		.OUT_PKT_BURST_TYPE_L          (40),
		.OUT_ST_DATA_W                 (64),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_006 (
		.clk                  (clk_clk),                                //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src10_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src10_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src10_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src10_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_006_src_data),             //          .data
		.out_channel          (width_adapter_006_src_channel),          //          .channel
		.out_valid            (width_adapter_006_src_valid),            //          .valid
		.out_ready            (width_adapter_006_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (24),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (33),
		.IN_PKT_BYTE_CNT_L             (31),
		.IN_PKT_TRANS_COMPRESSED_READ  (25),
		.IN_PKT_BURSTWRAP_H            (36),
		.IN_PKT_BURSTWRAP_L            (34),
		.IN_PKT_BURST_SIZE_H           (39),
		.IN_PKT_BURST_SIZE_L           (37),
		.IN_PKT_RESPONSE_STATUS_H      (63),
		.IN_PKT_RESPONSE_STATUS_L      (62),
		.IN_PKT_TRANS_EXCLUSIVE        (30),
		.IN_PKT_BURST_TYPE_H           (41),
		.IN_PKT_BURST_TYPE_L           (40),
		.IN_ST_DATA_W                  (64),
		.OUT_PKT_ADDR_H                (51),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (60),
		.OUT_PKT_BYTE_CNT_L            (58),
		.OUT_PKT_TRANS_COMPRESSED_READ (52),
		.OUT_PKT_BURST_SIZE_H          (66),
		.OUT_PKT_BURST_SIZE_L          (64),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (57),
		.OUT_PKT_BURST_TYPE_H          (68),
		.OUT_PKT_BURST_TYPE_L          (67),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_007 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_010_src_valid),             //      sink.valid
		.in_channel           (id_router_010_src_channel),           //          .channel
		.in_startofpacket     (id_router_010_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_010_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_010_src_ready),             //          .ready
		.in_data              (id_router_010_src_data),              //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_007_src_data),          //          .data
		.out_channel          (width_adapter_007_src_channel),       //          .channel
		.out_valid            (width_adapter_007_src_valid),         //          .valid
		.out_ready            (width_adapter_007_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	mysystem_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

endmodule
