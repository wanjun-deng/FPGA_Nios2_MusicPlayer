// mysystem.v

// Generated using ACDS version 13.1 162 at 2025.12.28.23:59:19

`timescale 1 ps / 1 ps
module mysystem (
		input  wire       clk_clk,                     //               clk.clk
		input  wire       reset_reset_n,               //             reset.reset_n
		output wire [7:0] led_export,                  //               led.export
		output wire       vib_export_export,           //        vib_export.export
		input  wire [3:0] keyboard_export_Row_i,       //   keyboard_export.Row_i
		output wire [3:0] keyboard_export_Col_o,       //                  .Col_o
		input  wire       ir_decode_export_iIR,        //  ir_decode_export.iIR
		output wire       ir_decode_export_Get_Flag_o, //                  .Get_Flag_o
		output wire       hex_driver_export_SH_CP,     // hex_driver_export.SH_CP
		output wire       hex_driver_export_ST_CP,     //                  .ST_CP
		output wire       hex_driver_export_DS         //                  .DS
	);

	wire   [7:0] mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_writedata;   // mm_interconnect_0:FreqSynth_IP_0_avalon_slave_0_writedata -> FreqSynth_IP_0:writedata
	wire   [1:0] mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_address;     // mm_interconnect_0:FreqSynth_IP_0_avalon_slave_0_address -> FreqSynth_IP_0:address
	wire         mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_chipselect;  // mm_interconnect_0:FreqSynth_IP_0_avalon_slave_0_chipselect -> FreqSynth_IP_0:chipselect
	wire         mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_write;       // mm_interconnect_0:FreqSynth_IP_0_avalon_slave_0_write -> FreqSynth_IP_0:write
	wire         mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_read;        // mm_interconnect_0:FreqSynth_IP_0_avalon_slave_0_read -> FreqSynth_IP_0:read
	wire   [7:0] mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_readdata;    // FreqSynth_IP_0:readdata -> mm_interconnect_0:FreqSynth_IP_0_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_keyboard_ip_0_avalon_slave_0_writedata;    // mm_interconnect_0:KeyBoard_IP_0_avalon_slave_0_writedata -> KeyBoard_IP_0:writedata
	wire   [0:0] mm_interconnect_0_keyboard_ip_0_avalon_slave_0_address;      // mm_interconnect_0:KeyBoard_IP_0_avalon_slave_0_address -> KeyBoard_IP_0:address
	wire         mm_interconnect_0_keyboard_ip_0_avalon_slave_0_chipselect;   // mm_interconnect_0:KeyBoard_IP_0_avalon_slave_0_chipselect -> KeyBoard_IP_0:chipselect
	wire         mm_interconnect_0_keyboard_ip_0_avalon_slave_0_write;        // mm_interconnect_0:KeyBoard_IP_0_avalon_slave_0_write -> KeyBoard_IP_0:write
	wire         mm_interconnect_0_keyboard_ip_0_avalon_slave_0_read;         // mm_interconnect_0:KeyBoard_IP_0_avalon_slave_0_read -> KeyBoard_IP_0:read
	wire   [7:0] mm_interconnect_0_keyboard_ip_0_avalon_slave_0_readdata;     // KeyBoard_IP_0:readdata -> mm_interconnect_0:KeyBoard_IP_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire         nios2_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [15:0] nios2_instruction_master_address;                            // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                               // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] nios2_instruction_master_readdata;                           // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_readdatavalid;                      // mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                      // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire   [2:0] mm_interconnect_0_pio_led_s1_address;                        // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_chipselect;                     // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire         mm_interconnect_0_pio_led_s1_write;                          // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                       // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire  [31:0] mm_interconnect_0_rom_s1_writedata;                          // mm_interconnect_0:rom_s1_writedata -> rom:writedata
	wire   [8:0] mm_interconnect_0_rom_s1_address;                            // mm_interconnect_0:rom_s1_address -> rom:address
	wire         mm_interconnect_0_rom_s1_chipselect;                         // mm_interconnect_0:rom_s1_chipselect -> rom:chipselect
	wire         mm_interconnect_0_rom_s1_clken;                              // mm_interconnect_0:rom_s1_clken -> rom:clken
	wire         mm_interconnect_0_rom_s1_write;                              // mm_interconnect_0:rom_s1_write -> rom:write
	wire  [31:0] mm_interconnect_0_rom_s1_readdata;                           // rom:readdata -> mm_interconnect_0:rom_s1_readdata
	wire         mm_interconnect_0_rom_s1_debugaccess;                        // mm_interconnect_0:rom_s1_debugaccess -> rom:debugaccess
	wire   [3:0] mm_interconnect_0_rom_s1_byteenable;                         // mm_interconnect_0:rom_s1_byteenable -> rom:byteenable
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                          // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                            // mm_interconnect_0:ram_s1_address -> ram:address
	wire         mm_interconnect_0_ram_s1_chipselect;                         // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire         mm_interconnect_0_ram_s1_clken;                              // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire         mm_interconnect_0_ram_s1_write;                              // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                           // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                         // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;               // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;              // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [7:0] mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_writedata;  // mm_interconnect_0:Hex_Driver_IP_0_avalon_slave_0_writedata -> Hex_Driver_IP_0:writedata
	wire   [2:0] mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_address;    // mm_interconnect_0:Hex_Driver_IP_0_avalon_slave_0_address -> Hex_Driver_IP_0:address
	wire         mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_chipselect; // mm_interconnect_0:Hex_Driver_IP_0_avalon_slave_0_chipselect -> Hex_Driver_IP_0:chipselect
	wire         mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_write;      // mm_interconnect_0:Hex_Driver_IP_0_avalon_slave_0_write -> Hex_Driver_IP_0:write
	wire         mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_read;       // mm_interconnect_0:Hex_Driver_IP_0_avalon_slave_0_read -> Hex_Driver_IP_0:read
	wire   [7:0] mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_readdata;   // Hex_Driver_IP_0:readdata -> mm_interconnect_0:Hex_Driver_IP_0_avalon_slave_0_readdata
	wire         nios2_data_master_waitrequest;                               // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire  [31:0] nios2_data_master_writedata;                                 // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [15:0] nios2_data_master_address;                                   // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire         nios2_data_master_write;                                     // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire         nios2_data_master_read;                                      // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire  [31:0] nios2_data_master_readdata;                                  // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_debugaccess;                               // nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire         nios2_data_master_readdatavalid;                             // mm_interconnect_0:nios2_data_master_readdatavalid -> nios2:d_readdatavalid
	wire   [3:0] nios2_data_master_byteenable;                                // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         mm_interconnect_0_nios2_jtag_debug_module_waitrequest;       // nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_writedata;         // mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_jtag_debug_module_address;           // mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_jtag_debug_module_write;             // mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_jtag_debug_module_read;              // mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_readdata;          // nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_debugaccess;       // mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_jtag_debug_module_byteenable;        // mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	wire   [7:0] mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_writedata;   // mm_interconnect_0:Ir_Decode_IP_0_avalon_slave_0_writedata -> Ir_Decode_IP_0:writedata
	wire   [2:0] mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_address;     // mm_interconnect_0:Ir_Decode_IP_0_avalon_slave_0_address -> Ir_Decode_IP_0:address
	wire         mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_chipselect;  // mm_interconnect_0:Ir_Decode_IP_0_avalon_slave_0_chipselect -> Ir_Decode_IP_0:chipselect
	wire         mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_write;       // mm_interconnect_0:Ir_Decode_IP_0_avalon_slave_0_write -> Ir_Decode_IP_0:write
	wire         mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_read;        // mm_interconnect_0:Ir_Decode_IP_0_avalon_slave_0_read -> Ir_Decode_IP_0:read
	wire   [7:0] mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_readdata;    // Ir_Decode_IP_0:readdata -> mm_interconnect_0:Ir_Decode_IP_0_avalon_slave_0_readdata
	wire         irq_mapper_receiver0_irq;                                    // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_d_irq_irq;                                             // irq_mapper:sender_irq -> nios2:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [FreqSynth_IP_0:reset_n, Hex_Driver_IP_0:reset_n, Ir_Decode_IP_0:reset_n, KeyBoard_IP_0:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_reset_n_reset_bridge_in_reset_reset, nios2:reset_n, pio_led:reset_n, ram:reset, rom:reset, rst_translator:in_reset, sysid:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2:reset_req, ram:reset_req, rom:reset_req, rst_translator:reset_req_in]
	wire         nios2_jtag_debug_module_reset_reset;                         // nios2:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	mysystem_nios2 nios2 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (nios2_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_data_master_read),                                //                          .read
		.d_readdata                            (nios2_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_data_master_write),                               //                          .write
		.d_writedata                           (nios2_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	mysystem_rom rom (
		.clk         (clk_clk),                              //   clk1.clk
		.address     (mm_interconnect_0_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_0_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req)    //       .reset_req
	);

	mysystem_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)   //       .reset_req
	);

	mysystem_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	mysystem_pio_led pio_led (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                               // external_connection.export
	);

	mysystem_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	mysystem_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	avalon_FreqSynth freqsynth_ip_0 (
		.clk        (clk_clk),                                                    //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                            //          reset.reset_n
		.address    (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_address),    // avalon_slave_0.address
		.writedata  (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_writedata),  //               .writedata
		.write      (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_write),      //               .write
		.read       (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_read),       //               .read
		.chipselect (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_chipselect), //               .chipselect
		.readdata   (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_readdata),   //               .readdata
		.vib        (vib_export_export)                                           //    conduit_end.export
	);

	avalon_KeyBoard keyboard_ip_0 (
		.clk             (clk_clk),                                                   //          clock.clk
		.reset_n         (~rst_controller_reset_out_reset),                           //          reset.reset_n
		.address         (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_address),    // avalon_slave_0.address
		.read            (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_read),       //               .read
		.chipselect      (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_chipselect), //               .chipselect
		.readdata        (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_readdata),   //               .readdata
		.writedata       (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_writedata),  //               .writedata
		.write           (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_write),      //               .write
		.Key_Board_Row_i (keyboard_export_Row_i),                                     //    conduit_end.export
		.Key_Board_Col_o (keyboard_export_Col_o)                                      //               .export
	);

	avalon_ir_decode ir_decode_ip_0 (
		.clk        (clk_clk),                                                    //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                            //          reset.reset_n
		.address    (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_address),    // avalon_slave_0.address
		.writedata  (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_writedata),  //               .writedata
		.write      (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_write),      //               .write
		.read       (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_read),       //               .read
		.chipselect (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_chipselect), //               .chipselect
		.readdata   (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_readdata),   //               .readdata
		.iIR        (ir_decode_export_iIR),                                       //    conduit_end.export
		.Get_Flag_o (ir_decode_export_Get_Flag_o)                                 //               .export
	);

	avalon_hex_top hex_driver_ip_0 (
		.clk        (clk_clk),                                                     //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                             //          reset.reset_n
		.address    (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_address),    // avalon_slave_0.address
		.writedata  (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_writedata),  //               .writedata
		.write      (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_write),      //               .write
		.read       (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_read),       //               .read
		.chipselect (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_chipselect), //               .chipselect
		.readdata   (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_readdata),   //               .readdata
		.SH_CP      (hex_driver_export_SH_CP),                                     //    conduit_end.export
		.ST_CP      (hex_driver_export_ST_CP),                                     //               .export
		.DS         (hex_driver_export_DS)                                         //               .export
	);

	mysystem_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                             (clk_clk),                                                     //                           clk_0_clk.clk
		.nios2_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_reset_n_reset_bridge_in_reset.reset
		.nios2_data_master_address                 (nios2_data_master_address),                                   //                   nios2_data_master.address
		.nios2_data_master_waitrequest             (nios2_data_master_waitrequest),                               //                                    .waitrequest
		.nios2_data_master_byteenable              (nios2_data_master_byteenable),                                //                                    .byteenable
		.nios2_data_master_read                    (nios2_data_master_read),                                      //                                    .read
		.nios2_data_master_readdata                (nios2_data_master_readdata),                                  //                                    .readdata
		.nios2_data_master_readdatavalid           (nios2_data_master_readdatavalid),                             //                                    .readdatavalid
		.nios2_data_master_write                   (nios2_data_master_write),                                     //                                    .write
		.nios2_data_master_writedata               (nios2_data_master_writedata),                                 //                                    .writedata
		.nios2_data_master_debugaccess             (nios2_data_master_debugaccess),                               //                                    .debugaccess
		.nios2_instruction_master_address          (nios2_instruction_master_address),                            //            nios2_instruction_master.address
		.nios2_instruction_master_waitrequest      (nios2_instruction_master_waitrequest),                        //                                    .waitrequest
		.nios2_instruction_master_read             (nios2_instruction_master_read),                               //                                    .read
		.nios2_instruction_master_readdata         (nios2_instruction_master_readdata),                           //                                    .readdata
		.nios2_instruction_master_readdatavalid    (nios2_instruction_master_readdatavalid),                      //                                    .readdatavalid
		.FreqSynth_IP_0_avalon_slave_0_address     (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_address),     //       FreqSynth_IP_0_avalon_slave_0.address
		.FreqSynth_IP_0_avalon_slave_0_write       (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_write),       //                                    .write
		.FreqSynth_IP_0_avalon_slave_0_read        (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_read),        //                                    .read
		.FreqSynth_IP_0_avalon_slave_0_readdata    (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_readdata),    //                                    .readdata
		.FreqSynth_IP_0_avalon_slave_0_writedata   (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_writedata),   //                                    .writedata
		.FreqSynth_IP_0_avalon_slave_0_chipselect  (mm_interconnect_0_freqsynth_ip_0_avalon_slave_0_chipselect),  //                                    .chipselect
		.Hex_Driver_IP_0_avalon_slave_0_address    (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_address),    //      Hex_Driver_IP_0_avalon_slave_0.address
		.Hex_Driver_IP_0_avalon_slave_0_write      (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_write),      //                                    .write
		.Hex_Driver_IP_0_avalon_slave_0_read       (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_read),       //                                    .read
		.Hex_Driver_IP_0_avalon_slave_0_readdata   (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_readdata),   //                                    .readdata
		.Hex_Driver_IP_0_avalon_slave_0_writedata  (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_writedata),  //                                    .writedata
		.Hex_Driver_IP_0_avalon_slave_0_chipselect (mm_interconnect_0_hex_driver_ip_0_avalon_slave_0_chipselect), //                                    .chipselect
		.Ir_Decode_IP_0_avalon_slave_0_address     (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_address),     //       Ir_Decode_IP_0_avalon_slave_0.address
		.Ir_Decode_IP_0_avalon_slave_0_write       (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_write),       //                                    .write
		.Ir_Decode_IP_0_avalon_slave_0_read        (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_read),        //                                    .read
		.Ir_Decode_IP_0_avalon_slave_0_readdata    (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_readdata),    //                                    .readdata
		.Ir_Decode_IP_0_avalon_slave_0_writedata   (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_writedata),   //                                    .writedata
		.Ir_Decode_IP_0_avalon_slave_0_chipselect  (mm_interconnect_0_ir_decode_ip_0_avalon_slave_0_chipselect),  //                                    .chipselect
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //       jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                    .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                    .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                    .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                    .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                    .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                    .chipselect
		.KeyBoard_IP_0_avalon_slave_0_address      (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_address),      //        KeyBoard_IP_0_avalon_slave_0.address
		.KeyBoard_IP_0_avalon_slave_0_write        (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_write),        //                                    .write
		.KeyBoard_IP_0_avalon_slave_0_read         (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_read),         //                                    .read
		.KeyBoard_IP_0_avalon_slave_0_readdata     (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_readdata),     //                                    .readdata
		.KeyBoard_IP_0_avalon_slave_0_writedata    (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_writedata),    //                                    .writedata
		.KeyBoard_IP_0_avalon_slave_0_chipselect   (mm_interconnect_0_keyboard_ip_0_avalon_slave_0_chipselect),   //                                    .chipselect
		.nios2_jtag_debug_module_address           (mm_interconnect_0_nios2_jtag_debug_module_address),           //             nios2_jtag_debug_module.address
		.nios2_jtag_debug_module_write             (mm_interconnect_0_nios2_jtag_debug_module_write),             //                                    .write
		.nios2_jtag_debug_module_read              (mm_interconnect_0_nios2_jtag_debug_module_read),              //                                    .read
		.nios2_jtag_debug_module_readdata          (mm_interconnect_0_nios2_jtag_debug_module_readdata),          //                                    .readdata
		.nios2_jtag_debug_module_writedata         (mm_interconnect_0_nios2_jtag_debug_module_writedata),         //                                    .writedata
		.nios2_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_jtag_debug_module_byteenable),        //                                    .byteenable
		.nios2_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_jtag_debug_module_waitrequest),       //                                    .waitrequest
		.nios2_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_jtag_debug_module_debugaccess),       //                                    .debugaccess
		.pio_led_s1_address                        (mm_interconnect_0_pio_led_s1_address),                        //                          pio_led_s1.address
		.pio_led_s1_write                          (mm_interconnect_0_pio_led_s1_write),                          //                                    .write
		.pio_led_s1_readdata                       (mm_interconnect_0_pio_led_s1_readdata),                       //                                    .readdata
		.pio_led_s1_writedata                      (mm_interconnect_0_pio_led_s1_writedata),                      //                                    .writedata
		.pio_led_s1_chipselect                     (mm_interconnect_0_pio_led_s1_chipselect),                     //                                    .chipselect
		.ram_s1_address                            (mm_interconnect_0_ram_s1_address),                            //                              ram_s1.address
		.ram_s1_write                              (mm_interconnect_0_ram_s1_write),                              //                                    .write
		.ram_s1_readdata                           (mm_interconnect_0_ram_s1_readdata),                           //                                    .readdata
		.ram_s1_writedata                          (mm_interconnect_0_ram_s1_writedata),                          //                                    .writedata
		.ram_s1_byteenable                         (mm_interconnect_0_ram_s1_byteenable),                         //                                    .byteenable
		.ram_s1_chipselect                         (mm_interconnect_0_ram_s1_chipselect),                         //                                    .chipselect
		.ram_s1_clken                              (mm_interconnect_0_ram_s1_clken),                              //                                    .clken
		.rom_s1_address                            (mm_interconnect_0_rom_s1_address),                            //                              rom_s1.address
		.rom_s1_write                              (mm_interconnect_0_rom_s1_write),                              //                                    .write
		.rom_s1_readdata                           (mm_interconnect_0_rom_s1_readdata),                           //                                    .readdata
		.rom_s1_writedata                          (mm_interconnect_0_rom_s1_writedata),                          //                                    .writedata
		.rom_s1_byteenable                         (mm_interconnect_0_rom_s1_byteenable),                         //                                    .byteenable
		.rom_s1_chipselect                         (mm_interconnect_0_rom_s1_chipselect),                         //                                    .chipselect
		.rom_s1_clken                              (mm_interconnect_0_rom_s1_clken),                              //                                    .clken
		.rom_s1_debugaccess                        (mm_interconnect_0_rom_s1_debugaccess),                        //                                    .debugaccess
		.sysid_control_slave_address               (mm_interconnect_0_sysid_control_slave_address),               //                 sysid_control_slave.address
		.sysid_control_slave_readdata              (mm_interconnect_0_sysid_control_slave_readdata),              //                                    .readdata
		.timer_0_s1_address                        (mm_interconnect_0_timer_0_s1_address),                        //                          timer_0_s1.address
		.timer_0_s1_write                          (mm_interconnect_0_timer_0_s1_write),                          //                                    .write
		.timer_0_s1_readdata                       (mm_interconnect_0_timer_0_s1_readdata),                       //                                    .readdata
		.timer_0_s1_writedata                      (mm_interconnect_0_timer_0_s1_writedata),                      //                                    .writedata
		.timer_0_s1_chipselect                     (mm_interconnect_0_timer_0_s1_chipselect)                      //                                    .chipselect
	);

	mysystem_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
