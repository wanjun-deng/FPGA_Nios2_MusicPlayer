// mysystem.v

// Generated using ACDS version 13.1 162 at 2025.12.26.12:21:06

`timescale 1 ps / 1 ps
module mysystem (
		input  wire        clk_clk,           //        clk.clk
		input  wire        reset_reset_n,     //      reset.reset_n
		output wire [7:0]  led_export,        //        led.export
		input  wire [7:0]  keyboard_export,   //   keyboard.export
		output wire [7:0]  onote_export,      //      onote.export
		output wire [7:0]  playing_export,    //    playing.export
		input  wire [15:0] irdata_export,     //     irdata.export
		input  wire [7:0]  irflag_export,     //     irflag.export
		output wire [7:0]  volumectrl_export, // volumectrl.export
		output wire [31:0] display_export     //    display.export
	);

	wire   [1:0] mm_interconnect_0_pio_irflag_s1_address;                     // mm_interconnect_0:pio_irflag_s1_address -> pio_irflag:address
	wire  [31:0] mm_interconnect_0_pio_irflag_s1_readdata;                    // pio_irflag:readdata -> mm_interconnect_0:pio_irflag_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_onote_s1_writedata;                    // mm_interconnect_0:pio_onote_s1_writedata -> pio_onote:writedata
	wire   [2:0] mm_interconnect_0_pio_onote_s1_address;                      // mm_interconnect_0:pio_onote_s1_address -> pio_onote:address
	wire         mm_interconnect_0_pio_onote_s1_chipselect;                   // mm_interconnect_0:pio_onote_s1_chipselect -> pio_onote:chipselect
	wire         mm_interconnect_0_pio_onote_s1_write;                        // mm_interconnect_0:pio_onote_s1_write -> pio_onote:write_n
	wire  [31:0] mm_interconnect_0_pio_onote_s1_readdata;                     // pio_onote:readdata -> mm_interconnect_0:pio_onote_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_volumectrl_s1_writedata;               // mm_interconnect_0:pio_volumectrl_s1_writedata -> pio_volumectrl:writedata
	wire   [2:0] mm_interconnect_0_pio_volumectrl_s1_address;                 // mm_interconnect_0:pio_volumectrl_s1_address -> pio_volumectrl:address
	wire         mm_interconnect_0_pio_volumectrl_s1_chipselect;              // mm_interconnect_0:pio_volumectrl_s1_chipselect -> pio_volumectrl:chipselect
	wire         mm_interconnect_0_pio_volumectrl_s1_write;                   // mm_interconnect_0:pio_volumectrl_s1_write -> pio_volumectrl:write_n
	wire  [31:0] mm_interconnect_0_pio_volumectrl_s1_readdata;                // pio_volumectrl:readdata -> mm_interconnect_0:pio_volumectrl_s1_readdata
	wire         nios2_data_master_waitrequest;                               // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire  [31:0] nios2_data_master_writedata;                                 // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [15:0] nios2_data_master_address;                                   // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire         nios2_data_master_write;                                     // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire         nios2_data_master_read;                                      // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire  [31:0] nios2_data_master_readdata;                                  // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_debugaccess;                               // nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire         nios2_data_master_readdatavalid;                             // mm_interconnect_0:nios2_data_master_readdatavalid -> nios2:d_readdatavalid
	wire   [3:0] nios2_data_master_byteenable;                                // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire  [31:0] mm_interconnect_0_pio_display_s1_writedata;                  // mm_interconnect_0:pio_display_s1_writedata -> pio_display:writedata
	wire   [2:0] mm_interconnect_0_pio_display_s1_address;                    // mm_interconnect_0:pio_display_s1_address -> pio_display:address
	wire         mm_interconnect_0_pio_display_s1_chipselect;                 // mm_interconnect_0:pio_display_s1_chipselect -> pio_display:chipselect
	wire         mm_interconnect_0_pio_display_s1_write;                      // mm_interconnect_0:pio_display_s1_write -> pio_display:write_n
	wire  [31:0] mm_interconnect_0_pio_display_s1_readdata;                   // pio_display:readdata -> mm_interconnect_0:pio_display_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_irdata_s1_address;                     // mm_interconnect_0:pio_irdata_s1_address -> pio_irdata:address
	wire  [31:0] mm_interconnect_0_pio_irdata_s1_readdata;                    // pio_irdata:readdata -> mm_interconnect_0:pio_irdata_s1_readdata
	wire  [31:0] mm_interconnect_0_rom_s1_writedata;                          // mm_interconnect_0:rom_s1_writedata -> rom:writedata
	wire   [8:0] mm_interconnect_0_rom_s1_address;                            // mm_interconnect_0:rom_s1_address -> rom:address
	wire         mm_interconnect_0_rom_s1_chipselect;                         // mm_interconnect_0:rom_s1_chipselect -> rom:chipselect
	wire         mm_interconnect_0_rom_s1_clken;                              // mm_interconnect_0:rom_s1_clken -> rom:clken
	wire         mm_interconnect_0_rom_s1_write;                              // mm_interconnect_0:rom_s1_write -> rom:write
	wire  [31:0] mm_interconnect_0_rom_s1_readdata;                           // rom:readdata -> mm_interconnect_0:rom_s1_readdata
	wire         mm_interconnect_0_rom_s1_debugaccess;                        // mm_interconnect_0:rom_s1_debugaccess -> rom:debugaccess
	wire   [3:0] mm_interconnect_0_rom_s1_byteenable;                         // mm_interconnect_0:rom_s1_byteenable -> rom:byteenable
	wire   [2:0] mm_interconnect_0_pio_keyboard_s1_address;                   // mm_interconnect_0:pio_keyboard_s1_address -> pio_keyboard:address
	wire  [31:0] mm_interconnect_0_pio_keyboard_s1_readdata;                  // pio_keyboard:readdata -> mm_interconnect_0:pio_keyboard_s1_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                      // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire   [2:0] mm_interconnect_0_pio_led_s1_address;                        // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_chipselect;                     // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire         mm_interconnect_0_pio_led_s1_write;                          // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                       // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire         nios2_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [15:0] nios2_instruction_master_address;                            // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                               // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] nios2_instruction_master_readdata;                           // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_readdatavalid;                      // mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	wire         mm_interconnect_0_nios2_jtag_debug_module_waitrequest;       // nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_writedata;         // mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_jtag_debug_module_address;           // mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_jtag_debug_module_write;             // mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_jtag_debug_module_read;              // mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_readdata;          // nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_debugaccess;       // mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_jtag_debug_module_byteenable;        // mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                          // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                            // mm_interconnect_0:ram_s1_address -> ram:address
	wire         mm_interconnect_0_ram_s1_chipselect;                         // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire         mm_interconnect_0_ram_s1_clken;                              // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire         mm_interconnect_0_ram_s1_write;                              // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                           // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                         // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_playing_s1_writedata;                  // mm_interconnect_0:pio_playing_s1_writedata -> pio_playing:writedata
	wire   [2:0] mm_interconnect_0_pio_playing_s1_address;                    // mm_interconnect_0:pio_playing_s1_address -> pio_playing:address
	wire         mm_interconnect_0_pio_playing_s1_chipselect;                 // mm_interconnect_0:pio_playing_s1_chipselect -> pio_playing:chipselect
	wire         mm_interconnect_0_pio_playing_s1_write;                      // mm_interconnect_0:pio_playing_s1_write -> pio_playing:write_n
	wire  [31:0] mm_interconnect_0_pio_playing_s1_readdata;                   // pio_playing:readdata -> mm_interconnect_0:pio_playing_s1_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;               // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;              // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire         irq_mapper_receiver0_irq;                                    // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_d_irq_irq;                                             // irq_mapper:sender_irq -> nios2:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_reset_n_reset_bridge_in_reset_reset, nios2:reset_n, pio_display:reset_n, pio_irdata:reset_n, pio_irflag:reset_n, pio_keyboard:reset_n, pio_led:reset_n, pio_onote:reset_n, pio_playing:reset_n, pio_volumectrl:reset_n, ram:reset, rom:reset, rst_translator:in_reset, sysid:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2:reset_req, ram:reset_req, rom:reset_req, rst_translator:reset_req_in]
	wire         nios2_jtag_debug_module_reset_reset;                         // nios2:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	mysystem_nios2 nios2 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (nios2_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_data_master_read),                                //                          .read
		.d_readdata                            (nios2_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_data_master_write),                               //                          .write
		.d_writedata                           (nios2_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	mysystem_rom rom (
		.clk         (clk_clk),                              //   clk1.clk
		.address     (mm_interconnect_0_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_0_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req)    //       .reset_req
	);

	mysystem_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)   //       .reset_req
	);

	mysystem_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	mysystem_pio_led pio_led (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                               // external_connection.export
	);

	mysystem_pio_keyboard pio_keyboard (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_pio_keyboard_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_keyboard_s1_readdata), //                    .readdata
		.in_port  (keyboard_export)                             // external_connection.export
	);

	mysystem_pio_onote pio_onote (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_onote_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_onote_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_onote_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_onote_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_onote_s1_readdata),   //                    .readdata
		.out_port   (onote_export)                               // external_connection.export
	);

	mysystem_pio_onote pio_playing (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pio_playing_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_playing_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_playing_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_playing_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_playing_s1_readdata),   //                    .readdata
		.out_port   (playing_export)                               // external_connection.export
	);

	mysystem_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	mysystem_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	mysystem_pio_irdata pio_irdata (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pio_irdata_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_irdata_s1_readdata), //                    .readdata
		.in_port  (irdata_export)                             // external_connection.export
	);

	mysystem_pio_irflag pio_irflag (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pio_irflag_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_irflag_s1_readdata), //                    .readdata
		.in_port  (irflag_export)                             // external_connection.export
	);

	mysystem_pio_onote pio_volumectrl (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_pio_volumectrl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_volumectrl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_volumectrl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_volumectrl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_volumectrl_s1_readdata),   //                    .readdata
		.out_port   (volumectrl_export)                               // external_connection.export
	);

	mysystem_pio_display pio_display (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pio_display_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_display_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_display_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_display_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_display_s1_readdata),   //                    .readdata
		.out_port   (display_export)                               // external_connection.export
	);

	mysystem_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                             (clk_clk),                                                     //                           clk_0_clk.clk
		.nios2_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_reset_n_reset_bridge_in_reset.reset
		.nios2_data_master_address                 (nios2_data_master_address),                                   //                   nios2_data_master.address
		.nios2_data_master_waitrequest             (nios2_data_master_waitrequest),                               //                                    .waitrequest
		.nios2_data_master_byteenable              (nios2_data_master_byteenable),                                //                                    .byteenable
		.nios2_data_master_read                    (nios2_data_master_read),                                      //                                    .read
		.nios2_data_master_readdata                (nios2_data_master_readdata),                                  //                                    .readdata
		.nios2_data_master_readdatavalid           (nios2_data_master_readdatavalid),                             //                                    .readdatavalid
		.nios2_data_master_write                   (nios2_data_master_write),                                     //                                    .write
		.nios2_data_master_writedata               (nios2_data_master_writedata),                                 //                                    .writedata
		.nios2_data_master_debugaccess             (nios2_data_master_debugaccess),                               //                                    .debugaccess
		.nios2_instruction_master_address          (nios2_instruction_master_address),                            //            nios2_instruction_master.address
		.nios2_instruction_master_waitrequest      (nios2_instruction_master_waitrequest),                        //                                    .waitrequest
		.nios2_instruction_master_read             (nios2_instruction_master_read),                               //                                    .read
		.nios2_instruction_master_readdata         (nios2_instruction_master_readdata),                           //                                    .readdata
		.nios2_instruction_master_readdatavalid    (nios2_instruction_master_readdatavalid),                      //                                    .readdatavalid
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //       jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                    .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                    .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                    .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                    .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                    .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                    .chipselect
		.nios2_jtag_debug_module_address           (mm_interconnect_0_nios2_jtag_debug_module_address),           //             nios2_jtag_debug_module.address
		.nios2_jtag_debug_module_write             (mm_interconnect_0_nios2_jtag_debug_module_write),             //                                    .write
		.nios2_jtag_debug_module_read              (mm_interconnect_0_nios2_jtag_debug_module_read),              //                                    .read
		.nios2_jtag_debug_module_readdata          (mm_interconnect_0_nios2_jtag_debug_module_readdata),          //                                    .readdata
		.nios2_jtag_debug_module_writedata         (mm_interconnect_0_nios2_jtag_debug_module_writedata),         //                                    .writedata
		.nios2_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_jtag_debug_module_byteenable),        //                                    .byteenable
		.nios2_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_jtag_debug_module_waitrequest),       //                                    .waitrequest
		.nios2_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_jtag_debug_module_debugaccess),       //                                    .debugaccess
		.pio_display_s1_address                    (mm_interconnect_0_pio_display_s1_address),                    //                      pio_display_s1.address
		.pio_display_s1_write                      (mm_interconnect_0_pio_display_s1_write),                      //                                    .write
		.pio_display_s1_readdata                   (mm_interconnect_0_pio_display_s1_readdata),                   //                                    .readdata
		.pio_display_s1_writedata                  (mm_interconnect_0_pio_display_s1_writedata),                  //                                    .writedata
		.pio_display_s1_chipselect                 (mm_interconnect_0_pio_display_s1_chipselect),                 //                                    .chipselect
		.pio_irdata_s1_address                     (mm_interconnect_0_pio_irdata_s1_address),                     //                       pio_irdata_s1.address
		.pio_irdata_s1_readdata                    (mm_interconnect_0_pio_irdata_s1_readdata),                    //                                    .readdata
		.pio_irflag_s1_address                     (mm_interconnect_0_pio_irflag_s1_address),                     //                       pio_irflag_s1.address
		.pio_irflag_s1_readdata                    (mm_interconnect_0_pio_irflag_s1_readdata),                    //                                    .readdata
		.pio_keyboard_s1_address                   (mm_interconnect_0_pio_keyboard_s1_address),                   //                     pio_keyboard_s1.address
		.pio_keyboard_s1_readdata                  (mm_interconnect_0_pio_keyboard_s1_readdata),                  //                                    .readdata
		.pio_led_s1_address                        (mm_interconnect_0_pio_led_s1_address),                        //                          pio_led_s1.address
		.pio_led_s1_write                          (mm_interconnect_0_pio_led_s1_write),                          //                                    .write
		.pio_led_s1_readdata                       (mm_interconnect_0_pio_led_s1_readdata),                       //                                    .readdata
		.pio_led_s1_writedata                      (mm_interconnect_0_pio_led_s1_writedata),                      //                                    .writedata
		.pio_led_s1_chipselect                     (mm_interconnect_0_pio_led_s1_chipselect),                     //                                    .chipselect
		.pio_onote_s1_address                      (mm_interconnect_0_pio_onote_s1_address),                      //                        pio_onote_s1.address
		.pio_onote_s1_write                        (mm_interconnect_0_pio_onote_s1_write),                        //                                    .write
		.pio_onote_s1_readdata                     (mm_interconnect_0_pio_onote_s1_readdata),                     //                                    .readdata
		.pio_onote_s1_writedata                    (mm_interconnect_0_pio_onote_s1_writedata),                    //                                    .writedata
		.pio_onote_s1_chipselect                   (mm_interconnect_0_pio_onote_s1_chipselect),                   //                                    .chipselect
		.pio_playing_s1_address                    (mm_interconnect_0_pio_playing_s1_address),                    //                      pio_playing_s1.address
		.pio_playing_s1_write                      (mm_interconnect_0_pio_playing_s1_write),                      //                                    .write
		.pio_playing_s1_readdata                   (mm_interconnect_0_pio_playing_s1_readdata),                   //                                    .readdata
		.pio_playing_s1_writedata                  (mm_interconnect_0_pio_playing_s1_writedata),                  //                                    .writedata
		.pio_playing_s1_chipselect                 (mm_interconnect_0_pio_playing_s1_chipselect),                 //                                    .chipselect
		.pio_volumectrl_s1_address                 (mm_interconnect_0_pio_volumectrl_s1_address),                 //                   pio_volumectrl_s1.address
		.pio_volumectrl_s1_write                   (mm_interconnect_0_pio_volumectrl_s1_write),                   //                                    .write
		.pio_volumectrl_s1_readdata                (mm_interconnect_0_pio_volumectrl_s1_readdata),                //                                    .readdata
		.pio_volumectrl_s1_writedata               (mm_interconnect_0_pio_volumectrl_s1_writedata),               //                                    .writedata
		.pio_volumectrl_s1_chipselect              (mm_interconnect_0_pio_volumectrl_s1_chipselect),              //                                    .chipselect
		.ram_s1_address                            (mm_interconnect_0_ram_s1_address),                            //                              ram_s1.address
		.ram_s1_write                              (mm_interconnect_0_ram_s1_write),                              //                                    .write
		.ram_s1_readdata                           (mm_interconnect_0_ram_s1_readdata),                           //                                    .readdata
		.ram_s1_writedata                          (mm_interconnect_0_ram_s1_writedata),                          //                                    .writedata
		.ram_s1_byteenable                         (mm_interconnect_0_ram_s1_byteenable),                         //                                    .byteenable
		.ram_s1_chipselect                         (mm_interconnect_0_ram_s1_chipselect),                         //                                    .chipselect
		.ram_s1_clken                              (mm_interconnect_0_ram_s1_clken),                              //                                    .clken
		.rom_s1_address                            (mm_interconnect_0_rom_s1_address),                            //                              rom_s1.address
		.rom_s1_write                              (mm_interconnect_0_rom_s1_write),                              //                                    .write
		.rom_s1_readdata                           (mm_interconnect_0_rom_s1_readdata),                           //                                    .readdata
		.rom_s1_writedata                          (mm_interconnect_0_rom_s1_writedata),                          //                                    .writedata
		.rom_s1_byteenable                         (mm_interconnect_0_rom_s1_byteenable),                         //                                    .byteenable
		.rom_s1_chipselect                         (mm_interconnect_0_rom_s1_chipselect),                         //                                    .chipselect
		.rom_s1_clken                              (mm_interconnect_0_rom_s1_clken),                              //                                    .clken
		.rom_s1_debugaccess                        (mm_interconnect_0_rom_s1_debugaccess),                        //                                    .debugaccess
		.sysid_control_slave_address               (mm_interconnect_0_sysid_control_slave_address),               //                 sysid_control_slave.address
		.sysid_control_slave_readdata              (mm_interconnect_0_sysid_control_slave_readdata),              //                                    .readdata
		.timer_0_s1_address                        (mm_interconnect_0_timer_0_s1_address),                        //                          timer_0_s1.address
		.timer_0_s1_write                          (mm_interconnect_0_timer_0_s1_write),                          //                                    .write
		.timer_0_s1_readdata                       (mm_interconnect_0_timer_0_s1_readdata),                       //                                    .readdata
		.timer_0_s1_writedata                      (mm_interconnect_0_timer_0_s1_writedata),                      //                                    .writedata
		.timer_0_s1_chipselect                     (mm_interconnect_0_timer_0_s1_chipselect)                      //                                    .chipselect
	);

	mysystem_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
